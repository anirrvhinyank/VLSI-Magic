magic
tech scmos
timestamp 1635336988
<< nwell >>
rect -8 -5 42 8
<< polysilicon >>
rect 1 6 4 8
rect 14 6 17 8
rect 32 6 35 8
rect 1 -9 4 -3
rect 14 -9 17 -3
rect 32 -9 35 -3
rect 2 -13 4 -9
rect 16 -13 17 -9
rect 26 -13 35 -9
rect 1 -28 4 -13
rect 14 -28 17 -13
rect 32 -28 35 -13
rect 1 -39 4 -37
rect 14 -39 17 -37
rect 32 -39 35 -37
<< ndiffusion >>
rect -6 -29 1 -28
rect -2 -33 1 -29
rect -6 -37 1 -33
rect 4 -29 14 -28
rect 4 -33 7 -29
rect 11 -33 14 -29
rect 4 -37 14 -33
rect 17 -29 22 -28
rect 17 -33 18 -29
rect 17 -37 22 -33
rect 27 -30 32 -28
rect 31 -34 32 -30
rect 27 -37 32 -34
rect 35 -30 40 -28
rect 35 -34 36 -30
rect 35 -37 40 -34
<< pdiffusion >>
rect -6 2 1 6
rect -6 -2 -5 2
rect -1 -2 1 2
rect -6 -3 1 -2
rect 4 -3 14 6
rect 17 4 23 6
rect 17 0 19 4
rect 17 -3 23 0
rect 27 4 32 6
rect 31 0 32 4
rect 27 -3 32 0
rect 35 4 40 6
rect 35 0 36 4
rect 35 -3 40 0
<< metal1 >>
rect -1 13 3 17
rect 7 13 11 17
rect 15 13 19 17
rect 23 13 27 17
rect -5 2 -1 13
rect 27 4 31 13
rect 19 -9 23 0
rect -8 -13 -2 -9
rect 7 -13 12 -9
rect 19 -13 22 -9
rect 36 -11 40 0
rect 19 -16 23 -13
rect 7 -20 23 -16
rect 36 -15 44 -11
rect 7 -29 11 -20
rect 36 -30 40 -15
rect -6 -44 -2 -33
rect 18 -44 22 -33
rect 27 -44 31 -34
rect -2 -48 2 -44
rect 6 -48 10 -44
rect 14 -48 18 -44
rect 22 -48 27 -44
<< ntransistor >>
rect 1 -37 4 -28
rect 14 -37 17 -28
rect 32 -37 35 -28
<< ptransistor >>
rect 1 -3 4 6
rect 14 -3 17 6
rect 32 -3 35 6
<< polycontact >>
rect -2 -13 2 -9
rect 12 -13 16 -9
rect 22 -13 26 -9
<< ndcontact >>
rect -6 -33 -2 -29
rect 7 -33 11 -29
rect 18 -33 22 -29
rect 27 -34 31 -30
rect 36 -34 40 -30
<< pdcontact >>
rect -5 -2 -1 2
rect 19 0 23 4
rect 27 0 31 4
rect 36 0 40 4
<< psubstratepcontact >>
rect -6 -48 -2 -44
rect 2 -48 6 -44
rect 10 -48 14 -44
rect 18 -48 22 -44
rect 27 -48 31 -44
<< nsubstratencontact >>
rect -5 13 -1 17
rect 3 13 7 17
rect 11 13 15 17
rect 19 13 23 17
rect 27 13 31 17
<< labels >>
rlabel metal1 -3 10 -3 10 3 Vdd
rlabel metal1 -5 -41 -5 -41 3 gnd
rlabel metal1 -5 -11 -5 -11 3 a
rlabel metal1 9 -11 9 -11 1 v
rlabel metal1 9 -11 9 -11 1 b
rlabel metal1 38 -12 38 -12 7 out2
<< end >>
