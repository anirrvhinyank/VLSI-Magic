* SPICE3 file created from inverterfile.ext - technology: scmos

.option scale=1u

M1000 vout vin gnd Gnd nfet w=9 l=3
+  ad=0 pd=0 as=0 ps=0
M1001 vout vin Vdd w_n8_n5# pfet w=9 l=3
+  ad=0 pd=0 as=0 ps=0
C0 gnd Gnd 3.38fF
C1 vout Gnd 5.08fF
C2 vin Gnd 9.96fF
C3 Vdd Gnd 2.63fF
