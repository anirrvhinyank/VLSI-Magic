magic
tech scmos
timestamp 1636226274
<< nwell >>
rect -21 1 1 11
rect 27 2 49 12
rect 62 -44 130 -34
rect 62 -109 130 -99
rect 62 -173 130 -163
rect 62 -245 130 -235
<< polysilicon >>
rect -11 9 -9 13
rect 37 10 39 14
rect -11 -13 -9 3
rect 37 -12 39 4
rect -11 -49 -9 -19
rect -11 -51 7 -49
rect 5 -179 7 -51
rect 37 -85 39 -18
rect 72 -36 74 -32
rect 86 -36 88 -6
rect 118 -36 120 -32
rect 72 -58 74 -42
rect 86 -58 88 -42
rect 118 -49 120 -42
rect 117 -53 120 -49
rect 118 -58 120 -53
rect 72 -66 74 -64
rect 86 -80 88 -64
rect 118 -66 120 -64
rect 86 -82 164 -80
rect 37 -87 88 -85
rect 37 -89 39 -87
rect 36 -91 40 -89
rect 72 -101 74 -99
rect 86 -101 88 -87
rect 162 -90 164 -82
rect 118 -101 120 -99
rect 72 -123 74 -107
rect 86 -123 88 -107
rect 118 -114 120 -107
rect 117 -118 120 -114
rect 118 -123 120 -118
rect 72 -131 74 -129
rect 86 -131 88 -129
rect 118 -131 120 -129
rect 162 -142 164 -94
rect 86 -144 164 -142
rect 72 -165 74 -163
rect 86 -165 88 -144
rect 118 -165 120 -163
rect 72 -179 74 -171
rect 5 -183 21 -179
rect 52 -183 74 -179
rect 5 -251 7 -183
rect 72 -187 74 -183
rect 86 -187 88 -171
rect 118 -178 120 -171
rect 117 -182 120 -178
rect 118 -187 120 -182
rect 72 -195 74 -193
rect 86 -195 88 -193
rect 118 -195 120 -193
rect 72 -237 74 -235
rect 86 -237 88 -219
rect 118 -237 120 -235
rect 72 -251 74 -243
rect 5 -253 74 -251
rect 72 -259 74 -253
rect 86 -259 88 -243
rect 118 -250 120 -243
rect 117 -254 120 -250
rect 118 -259 120 -254
rect 72 -267 74 -265
rect 86 -267 88 -265
rect 118 -267 120 -265
<< ndiffusion >>
rect 29 -13 37 -12
rect -19 -14 -11 -13
rect -15 -18 -11 -14
rect -19 -19 -11 -18
rect -9 -14 -1 -13
rect -9 -18 -5 -14
rect 33 -17 37 -13
rect 29 -18 37 -17
rect 39 -13 47 -12
rect 39 -17 43 -13
rect 39 -18 47 -17
rect -9 -19 -1 -18
rect 64 -59 72 -58
rect 68 -63 72 -59
rect 64 -64 72 -63
rect 74 -64 86 -58
rect 88 -59 96 -58
rect 88 -63 92 -59
rect 88 -64 96 -63
rect 110 -59 118 -58
rect 114 -63 118 -59
rect 110 -64 118 -63
rect 120 -59 128 -58
rect 120 -63 124 -59
rect 120 -64 128 -63
rect 64 -124 72 -123
rect 68 -128 72 -124
rect 64 -129 72 -128
rect 74 -129 86 -123
rect 88 -124 96 -123
rect 88 -128 92 -124
rect 88 -129 96 -128
rect 110 -124 118 -123
rect 114 -128 118 -124
rect 110 -129 118 -128
rect 120 -124 128 -123
rect 120 -128 124 -124
rect 120 -129 128 -128
rect 64 -188 72 -187
rect 68 -192 72 -188
rect 64 -193 72 -192
rect 74 -193 86 -187
rect 88 -188 96 -187
rect 88 -192 92 -188
rect 88 -193 96 -192
rect 110 -188 118 -187
rect 114 -192 118 -188
rect 110 -193 118 -192
rect 120 -188 128 -187
rect 120 -192 124 -188
rect 120 -193 128 -192
rect 64 -260 72 -259
rect 68 -264 72 -260
rect 64 -265 72 -264
rect 74 -265 86 -259
rect 88 -260 96 -259
rect 88 -264 92 -260
rect 88 -265 96 -264
rect 110 -260 118 -259
rect 114 -264 118 -260
rect 110 -265 118 -264
rect 120 -260 128 -259
rect 120 -264 124 -260
rect 120 -265 128 -264
<< pdiffusion >>
rect 29 9 37 10
rect -19 8 -11 9
rect -15 4 -11 8
rect -19 3 -11 4
rect -9 8 -1 9
rect -9 4 -5 8
rect 33 5 37 9
rect 29 4 37 5
rect 39 9 47 10
rect 39 5 43 9
rect 39 4 47 5
rect -9 3 -1 4
rect 64 -37 72 -36
rect 68 -41 72 -37
rect 64 -42 72 -41
rect 74 -37 86 -36
rect 74 -41 78 -37
rect 82 -41 86 -37
rect 74 -42 86 -41
rect 88 -37 96 -36
rect 88 -41 92 -37
rect 88 -42 96 -41
rect 110 -37 118 -36
rect 114 -41 118 -37
rect 110 -42 118 -41
rect 120 -37 128 -36
rect 120 -41 124 -37
rect 120 -42 128 -41
rect 64 -102 72 -101
rect 68 -106 72 -102
rect 64 -107 72 -106
rect 74 -102 86 -101
rect 74 -106 78 -102
rect 82 -106 86 -102
rect 74 -107 86 -106
rect 88 -102 96 -101
rect 88 -106 92 -102
rect 88 -107 96 -106
rect 110 -102 118 -101
rect 114 -106 118 -102
rect 110 -107 118 -106
rect 120 -102 128 -101
rect 120 -106 124 -102
rect 120 -107 128 -106
rect 64 -166 72 -165
rect 68 -170 72 -166
rect 64 -171 72 -170
rect 74 -166 86 -165
rect 74 -170 78 -166
rect 82 -170 86 -166
rect 74 -171 86 -170
rect 88 -166 96 -165
rect 88 -170 92 -166
rect 88 -171 96 -170
rect 110 -166 118 -165
rect 114 -170 118 -166
rect 110 -171 118 -170
rect 120 -166 128 -165
rect 120 -170 124 -166
rect 120 -171 128 -170
rect 64 -238 72 -237
rect 68 -242 72 -238
rect 64 -243 72 -242
rect 74 -238 86 -237
rect 74 -242 78 -238
rect 82 -242 86 -238
rect 74 -243 86 -242
rect 88 -238 96 -237
rect 88 -242 92 -238
rect 88 -243 96 -242
rect 110 -238 118 -237
rect 114 -242 118 -238
rect 110 -243 118 -242
rect 120 -238 128 -237
rect 120 -242 124 -238
rect 120 -243 128 -242
<< metal1 >>
rect -27 18 191 22
rect -19 8 -15 18
rect 29 9 33 18
rect -5 -3 -1 4
rect 43 -2 47 5
rect -5 -7 23 -3
rect -5 -14 -1 -7
rect -19 -23 -15 -18
rect -27 -27 -18 -23
rect -1 -27 11 -23
rect -27 -70 -23 -27
rect 19 -49 23 -7
rect 43 -6 84 -2
rect 43 -13 47 -6
rect 29 -23 33 -17
rect 31 -27 33 -23
rect 187 -26 191 18
rect 64 -30 191 -26
rect 64 -37 68 -30
rect 110 -37 114 -30
rect 78 -49 82 -41
rect 124 -49 128 -41
rect 19 -53 68 -49
rect 78 -53 113 -49
rect 124 -53 134 -49
rect -27 -74 9 -70
rect -27 -133 -23 -74
rect 19 -114 23 -53
rect 92 -59 96 -53
rect 124 -59 128 -53
rect 64 -70 68 -63
rect 110 -70 114 -63
rect 33 -74 114 -70
rect 187 -90 191 -30
rect 36 -101 40 -95
rect 64 -94 191 -90
rect 64 -102 68 -94
rect 92 -102 96 -94
rect 110 -102 114 -94
rect 78 -114 82 -106
rect 124 -114 128 -106
rect 19 -118 68 -114
rect 78 -118 113 -114
rect 124 -118 134 -114
rect 92 -124 96 -118
rect 124 -124 128 -118
rect 64 -133 68 -128
rect 110 -133 114 -128
rect -27 -137 114 -133
rect -27 -197 -23 -137
rect 187 -150 191 -94
rect 64 -154 191 -150
rect 64 -166 68 -154
rect 92 -166 96 -154
rect 110 -166 114 -154
rect 78 -178 82 -170
rect 124 -178 128 -170
rect 25 -183 48 -179
rect 78 -182 113 -178
rect 124 -182 134 -178
rect 92 -188 96 -182
rect 124 -188 128 -182
rect 64 -197 68 -192
rect 110 -197 114 -192
rect -27 -201 114 -197
rect -27 -281 -23 -201
rect 85 -215 89 -208
rect 187 -223 191 -154
rect 64 -227 191 -223
rect 64 -238 68 -227
rect 92 -238 96 -227
rect 110 -238 114 -227
rect 78 -250 82 -242
rect 124 -250 128 -242
rect 78 -254 113 -250
rect 124 -254 134 -250
rect 92 -260 96 -254
rect 124 -260 128 -254
rect 64 -281 68 -264
rect 110 -281 114 -264
rect -27 -285 114 -281
<< metal2 >>
rect -14 -27 -5 -23
rect 15 -27 27 -23
rect 13 -74 29 -70
rect 36 -204 40 -105
rect 36 -208 85 -204
<< ntransistor >>
rect -11 -19 -9 -13
rect 37 -18 39 -12
rect 72 -64 74 -58
rect 86 -64 88 -58
rect 118 -64 120 -58
rect 72 -129 74 -123
rect 86 -129 88 -123
rect 118 -129 120 -123
rect 72 -193 74 -187
rect 86 -193 88 -187
rect 118 -193 120 -187
rect 72 -265 74 -259
rect 86 -265 88 -259
rect 118 -265 120 -259
<< ptransistor >>
rect -11 3 -9 9
rect 37 4 39 10
rect 72 -42 74 -36
rect 86 -42 88 -36
rect 118 -42 120 -36
rect 72 -107 74 -101
rect 86 -107 88 -101
rect 118 -107 120 -101
rect 72 -171 74 -165
rect 86 -171 88 -165
rect 118 -171 120 -165
rect 72 -243 74 -237
rect 86 -243 88 -237
rect 118 -243 120 -237
<< polycontact >>
rect 84 -6 88 -2
rect 68 -53 72 -49
rect 113 -53 117 -49
rect 36 -95 40 -91
rect 68 -118 72 -114
rect 113 -118 117 -114
rect 21 -183 25 -179
rect 48 -183 52 -179
rect 113 -182 117 -178
rect 85 -219 89 -215
rect 113 -254 117 -250
<< ndcontact >>
rect -19 -18 -15 -14
rect -5 -18 -1 -14
rect 29 -17 33 -13
rect 43 -17 47 -13
rect 64 -63 68 -59
rect 92 -63 96 -59
rect 110 -63 114 -59
rect 124 -63 128 -59
rect 64 -128 68 -124
rect 92 -128 96 -124
rect 110 -128 114 -124
rect 124 -128 128 -124
rect 64 -192 68 -188
rect 92 -192 96 -188
rect 110 -192 114 -188
rect 124 -192 128 -188
rect 64 -264 68 -260
rect 92 -264 96 -260
rect 110 -264 114 -260
rect 124 -264 128 -260
<< pdcontact >>
rect -19 4 -15 8
rect -5 4 -1 8
rect 29 5 33 9
rect 43 5 47 9
rect 64 -41 68 -37
rect 78 -41 82 -37
rect 92 -41 96 -37
rect 110 -41 114 -37
rect 124 -41 128 -37
rect 64 -106 68 -102
rect 78 -106 82 -102
rect 92 -106 96 -102
rect 110 -106 114 -102
rect 124 -106 128 -102
rect 64 -170 68 -166
rect 78 -170 82 -166
rect 92 -170 96 -166
rect 110 -170 114 -166
rect 124 -170 128 -166
rect 64 -242 68 -238
rect 78 -242 82 -238
rect 92 -242 96 -238
rect 110 -242 114 -238
rect 124 -242 128 -238
<< m2contact >>
rect -18 -27 -14 -23
rect -5 -27 -1 -23
rect 11 -27 15 -23
rect 27 -27 31 -23
rect 9 -74 13 -70
rect 29 -74 33 -70
rect 36 -105 40 -101
rect 85 -208 89 -204
<< labels >>
rlabel metal1 -17 20 -17 20 5 vdd
rlabel polysilicon 38 13 38 13 1 a0
rlabel metal1 132 -51 132 -51 1 d0
rlabel metal1 131 -116 131 -116 1 d1
rlabel metal1 132 -180 132 -180 1 d2
rlabel metal1 130 -252 130 -252 1 d3
rlabel metal1 73 -4 73 -4 1 a0'
rlabel metal1 10 -282 10 -282 1 gnd
rlabel metal1 22 -50 22 -50 1 a1'
rlabel polysilicon -10 12 -10 12 1 a1
<< end >>
