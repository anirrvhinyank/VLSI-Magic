magic
tech scmos
timestamp 1635355844
<< nwell >>
rect -60 1 26 14
<< polysilicon >>
rect -65 25 -28 27
rect -65 -37 -63 25
rect -53 12 -51 14
rect -30 12 -28 25
rect -6 12 -4 14
rect 17 12 19 14
rect -53 -16 -51 3
rect -30 -1 -28 3
rect -6 -9 -4 3
rect 17 -9 19 3
rect -10 -13 -4 -9
rect 12 -13 19 -9
rect 35 -13 42 -9
rect -53 -18 -28 -16
rect -53 -24 -51 -22
rect -30 -24 -28 -18
rect -6 -24 -4 -13
rect 17 -24 19 -13
rect -53 -37 -51 -33
rect -65 -39 -51 -37
rect -53 -52 -51 -39
rect -30 -46 -28 -33
rect -6 -35 -4 -33
rect 17 -46 19 -33
rect -30 -48 19 -46
rect 40 -52 42 -13
rect -53 -54 42 -52
<< ndiffusion >>
rect -58 -27 -53 -24
rect -54 -31 -53 -27
rect -58 -33 -53 -31
rect -51 -27 -46 -24
rect -51 -31 -50 -27
rect -51 -33 -46 -31
rect -35 -27 -30 -24
rect -31 -31 -30 -27
rect -35 -33 -30 -31
rect -28 -27 -23 -24
rect -28 -31 -27 -27
rect -28 -33 -23 -31
rect -11 -27 -6 -24
rect -7 -31 -6 -27
rect -11 -33 -6 -31
rect -4 -27 1 -24
rect -4 -31 -3 -27
rect -4 -33 1 -31
rect 12 -27 17 -24
rect 16 -31 17 -27
rect 12 -33 17 -31
rect 19 -27 24 -24
rect 19 -31 20 -27
rect 19 -33 24 -31
<< pdiffusion >>
rect -58 10 -53 12
rect -54 6 -53 10
rect -58 3 -53 6
rect -51 10 -46 12
rect -51 6 -50 10
rect -51 3 -46 6
rect -35 10 -30 12
rect -31 6 -30 10
rect -35 3 -30 6
rect -28 10 -23 12
rect -28 6 -27 10
rect -28 3 -23 6
rect -11 10 -6 12
rect -7 6 -6 10
rect -11 3 -6 6
rect -4 10 1 12
rect -4 6 -3 10
rect -4 3 1 6
rect 12 10 17 12
rect 16 6 17 10
rect 12 3 17 6
rect 19 10 24 12
rect 19 6 20 10
rect 19 3 24 6
<< metal1 >>
rect -58 30 -15 34
rect -58 10 -54 30
rect -58 -27 -54 6
rect -58 -32 -54 -31
rect -50 17 -23 21
rect -50 10 -46 17
rect -50 -27 -46 6
rect -50 -32 -46 -31
rect -35 10 -31 11
rect -35 -27 -31 6
rect -35 -39 -31 -31
rect -27 10 -23 17
rect -27 -27 -23 6
rect -19 -9 -15 30
rect -11 20 16 24
rect -11 10 -7 20
rect -3 10 1 11
rect 12 10 16 20
rect 20 10 24 11
rect -19 -13 -14 -9
rect -3 -16 1 6
rect -27 -32 -23 -31
rect -18 -20 1 -16
rect -18 -39 -14 -20
rect -3 -27 1 -20
rect 20 -9 24 6
rect 20 -13 31 -9
rect 20 -27 24 -13
rect -35 -43 -14 -39
rect -11 -41 -7 -31
rect -3 -32 1 -31
rect 12 -41 16 -31
rect 20 -32 24 -31
rect -11 -45 16 -41
<< ntransistor >>
rect -53 -33 -51 -24
rect -30 -33 -28 -24
rect -6 -33 -4 -24
rect 17 -33 19 -24
<< ptransistor >>
rect -53 3 -51 12
rect -30 3 -28 12
rect -6 3 -4 12
rect 17 3 19 12
<< polycontact >>
rect -14 -13 -10 -9
rect 31 -13 35 -9
<< ndcontact >>
rect -58 -31 -54 -27
rect -50 -31 -46 -27
rect -35 -31 -31 -27
rect -27 -31 -23 -27
rect -11 -31 -7 -27
rect -3 -31 1 -27
rect 12 -31 16 -27
rect 20 -31 24 -27
<< pdcontact >>
rect -58 6 -54 10
rect -50 6 -46 10
rect -35 6 -31 10
rect -27 6 -23 10
rect -11 6 -7 10
rect -3 6 1 10
rect 12 6 16 10
rect 20 6 24 10
<< labels >>
rlabel polycontact -12 -11 -12 -11 1 va
rlabel metal1 -1 -11 -1 -11 1 vai
rlabel polysilicon 15 -11 15 -11 1 vb
rlabel polycontact 33 -11 33 -11 1 vbi
rlabel metal1 3 -43 3 -43 1 gnd
rlabel metal1 -38 19 -38 19 1 vout
rlabel metal1 2 22 2 22 1 vdd
<< end >>
