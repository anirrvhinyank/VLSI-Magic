* SPICE3 file created from fulladder4hope.ext - technology: scmos

.option scale=1u

M1000 a_414_38# a_268_108# a_414_72# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1001 a_n76_106# a_n266_146# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1002 a_78_n140# a_n118_n144# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1003 vdd cin a_78_148# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1004 a_218_n42# a_78_n6# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1005 vdd b2 a_717_148# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1006 a_1061_150# a_865_n142# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1007 a_907_108# a_717_148# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 a_717_n40# a2 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 vdd a_1575_46# a_2083_n2# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 a_1061_n138# a_865_n142# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1011 a_1739_n104# a3 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1012 a_3066_0# a_2870_n138# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1013 a_n266_n108# a1 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1014 gnd a_1879_n40# a_1887_n140# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1015 a_1397_40# a_1251_110# a_1397_74# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 a_1739_150# a3 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1017 a_78_n140# cin a_78_n106# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1018 a_2722_n102# a4 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1019 gnd b2 a_717_n140# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1020 a_907_108# a_717_148# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1021 gnd a_2862_n38# a_2870_n138# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1022 a_78_n40# a_n118_n144# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1023 a_226_n108# a_78_n140# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1024 vdd a_592_44# a_1061_150# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1025 a_2083_n36# a_1887_n140# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1026 a_2083_n136# a_1887_n140# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1027 a_2273_112# a_2083_152# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1028 a_717_148# a2 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1029 a_1879_n40# a_1739_n4# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1030 gnd a_3256_114# a_3402_44# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1031 a_414_72# a_n76_106# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1032 vdd b3 a_1739_150# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1033 gnd a_592_44# a_1061_n138# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1034 a_1739_n138# b3 a_1739_n104# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1035 a_n118_n110# a_n266_n142# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1036 a_2912_112# a_2722_152# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1037 a_n76_106# a_n266_146# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1038 gnd a_268_108# a_414_38# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1039 a_1061_n38# a_865_n142# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 a_857_n42# a_717_n6# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1041 a_3066_n34# a_2870_n138# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1042 s2 a_1061_n138# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1043 cout a_3402_44# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1044 vdd b4 a_2722_n2# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1045 s2 a_1201_n40# a_1209_n106# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1046 a_2597_48# a_2419_42# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1047 a_1201_n40# a_1061_n4# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1048 gnd a_218_n42# s1 Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1049 a_1061_116# a_865_n142# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1050 a_3214_n102# a_3066_n134# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1051 a_2722_n2# b4 a_2722_n36# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1052 a_2083_n2# a_1575_46# a_2083_n36# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1053 a_78_148# a_n118_n144# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1054 a_592_44# a_414_38# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1055 a_717_n106# a2 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1056 gnd a_2273_112# a_2419_42# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1057 a_3066_120# a_2870_n138# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1058 a_1739_n38# a3 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1059 a_2083_152# a_1887_n140# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1060 gnd a_1575_46# a_2083_n136# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1061 a_1739_116# a3 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1062 a_2597_48# a_2419_42# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1063 a_1397_40# a_907_108# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1064 a_1061_n4# a_592_44# a_1061_n38# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1065 a_3066_0# a_2597_48# a_3066_n34# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1066 gnd a_857_n42# a_865_n142# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1067 a_n266_n42# a1 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1068 a_n126_n44# a_n266_n8# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1069 a_1575_46# a_1397_40# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1070 s3 a_2083_n136# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1071 a_1739_n4# a3 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1072 s3 a_2223_n38# a_2231_n104# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1073 a_n266_112# a1 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1074 a_1061_150# a_592_44# a_1061_116# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1075 a_3402_78# a_2912_112# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1076 a_3066_154# a_2597_48# a_3066_120# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1077 a_1739_n4# b3 a_1739_n38# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1078 a_3256_114# a_3066_154# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1079 a_2722_n36# a4 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1080 a_717_n6# a2 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1081 vdd a_1575_46# a_2083_152# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1082 vdd b4 a_2722_152# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1083 s4 a_3206_n36# a_3214_n102# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1084 a_2912_112# a_2722_152# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1085 a_2419_76# a_1929_110# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1086 a_1739_150# b3 a_1739_116# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1087 a_1061_n4# a_865_n142# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1088 a_414_38# a_n76_106# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1089 a_1739_n138# a3 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1090 a_865_n142# a_717_n140# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1091 cout a_3402_44# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1092 a_3066_n100# a_2870_n138# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1093 a_n266_n8# b1 a_n266_n42# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1094 a_3066_n134# a_2870_n138# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1095 a_592_44# a_414_38# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1096 a_n266_146# b1 a_n266_112# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1097 a_1887_n106# a_1739_n138# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1098 a_2722_n136# a4 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1099 gnd cin a_78_n140# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1100 a_2722_n136# b4 a_2722_n102# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1101 a_78_n6# a_n118_n144# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1102 vdd cin a_78_n6# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1103 a_2223_n38# a_2083_n2# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1104 a_2083_118# a_1887_n140# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1105 a_2870_n104# a_2722_n136# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1106 s1 a_218_n42# a_226_n108# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1107 a_78_148# cin a_78_114# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1108 a_717_148# b2 a_717_114# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1109 a_3066_n134# a_2597_48# a_3066_n100# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1110 a_1575_46# a_1397_40# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1111 a_2722_152# a4 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 gnd a_n126_n44# a_n118_n144# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1113 a_1201_n40# a_1061_n4# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1114 a_n266_n8# a1 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1115 a_78_n106# a_n118_n144# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1116 gnd b1 a_n266_n142# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1117 gnd b3 a_1739_n138# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1118 a_3256_114# a_3066_154# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1119 gnd a_1251_110# a_1397_40# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1120 a_3206_n36# a_3066_0# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1121 a_1061_n104# a_865_n142# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1122 a_n126_n44# a_n266_n8# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1123 vdd b3 a_1739_n4# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1124 gnd a_2597_48# a_3066_n134# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1125 a_865_n142# a_857_n42# a_865_n108# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1126 a_1879_n40# a_1739_n4# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1127 gnd a_1201_n40# s2 Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1128 a_1887_n140# a_1879_n40# a_1887_n106# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1129 a_2083_152# a_1575_46# a_2083_118# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 a_3402_44# a_3256_114# a_3402_78# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1131 a_2722_152# b4 a_2722_118# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1132 a_1251_110# a_1061_150# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1133 a_218_n42# a_78_n6# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1134 s4 a_3066_n134# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1135 a_857_n42# a_717_n6# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1136 a_717_n140# a2 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1137 a_717_n140# b2 a_717_n106# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1138 a_717_114# a2 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1139 vdd a_592_44# a_1061_n4# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1140 a_2870_n138# a_2862_n38# a_2870_n104# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1141 a_1929_110# a_1739_150# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1142 a_2862_n38# a_2722_n2# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1143 a_865_n108# a_717_n140# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1144 vdd b2 a_717_n6# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1145 a_2419_42# a_2273_112# a_2419_76# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1146 a_2083_n102# a_1887_n140# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1147 a_2083_n2# a_1887_n140# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1148 a_n266_n142# a1 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1149 a_3066_154# a_2870_n138# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1150 a_2223_n38# a_2083_n2# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1151 a_268_108# a_78_148# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1152 gnd a_2223_n38# s3 Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1153 a_2862_n38# a_2722_n2# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1154 a_1397_74# a_907_108# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1155 a_1061_n138# a_592_44# a_1061_n104# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1156 vdd b1 a_n266_n8# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1157 a_78_114# a_n118_n144# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1158 a_2722_118# a4 gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1159 a_1209_n106# a_1061_n138# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1160 gnd a_3206_n36# s4 Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1161 s1 a_78_n140# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1162 a_n266_146# a1 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1163 a_3206_n36# a_3066_0# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1164 a_268_108# a_78_148# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1165 vdd a_2597_48# a_3066_154# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1166 a_78_n6# cin a_78_n40# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1167 a_n118_n144# a_n126_n44# a_n118_n110# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1168 a_717_n6# b2 a_717_n40# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1169 a_1251_110# a_1061_150# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1170 a_n266_n142# b1 a_n266_n108# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1171 a_1887_n140# a_1739_n138# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1172 a_2083_n136# a_1575_46# a_2083_n102# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1173 a_3402_44# a_2912_112# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1174 gnd b4 a_2722_n136# Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1175 a_2722_n2# a4 vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1176 a_n118_n144# a_n266_n142# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1177 a_1929_110# a_1739_150# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1178 a_2231_n104# a_2083_n136# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1179 vdd a_2597_48# a_3066_0# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1180 a_2273_112# a_2083_152# vdd Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1181 vdd b1 a_n266_146# Vdd pfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1182 a_2870_n138# a_2722_n136# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1183 a_2419_42# a_1929_110# gnd Gnd nfet w=10 l=4
+  ad=0 pd=0 as=0 ps=0
C0 a_268_108# gnd 5.70fF
C1 a_268_108# m2_472_6# 4.50fF
C2 a_2273_112# m2_2477_10# 4.50fF
C3 a1 vdd 3.60fF
C4 vdd a3 3.60fF
C5 vdd a_865_n142# 3.60fF
C6 cin vdd 3.60fF
C7 vdd a_1929_110# 11.22fF
C8 vdd a_3256_114# 12.36fF
C9 a_n118_n144# vdd 3.60fF
C10 vdd a_1887_n140# 3.60fF
C11 gnd b4 3.60fF
C12 gnd a2 3.60fF
C13 vdd a_907_108# 11.22fF
C14 a1 gnd 3.60fF
C15 gnd a3 3.60fF
C16 gnd a_865_n142# 4.80fF
C17 vdd a_2597_48# 4.80fF
C18 cin gnd 3.60fF
C19 gnd a_3256_114# 5.70fF
C20 a_n118_n144# gnd 4.80fF
C21 gnd a_1887_n140# 4.80fF
C22 a_592_44# vdd 4.80fF
C23 vdd a4 3.60fF
C24 gnd a_2597_48# 3.60fF
C25 a_1251_110# m2_1455_8# 4.50fF
C26 vdd a_2912_112# 10.02fF
C27 vdd a_2870_n138# 3.60fF
C28 vdd b2 3.60fF
C29 a_592_44# gnd 3.60fF
C30 b1 vdd 3.60fF
C31 vdd b3 3.60fF
C32 gnd a4 3.60fF
C33 vdd a_1575_46# 4.80fF
C34 a_n76_106# vdd 11.22fF
C35 gnd a_2870_n138# 4.80fF
C36 gnd b2 3.60fF
C37 vdd a_2273_112# 12.36fF
C38 b1 gnd 3.60fF
C39 gnd b3 3.60fF
C40 gnd a_1575_46# 3.60fF
C41 vdd a_1251_110# 12.36fF
C42 vdd a_268_108# 12.36fF
C43 gnd a_2273_112# 5.70fF
C44 a_3256_114# m2_3460_12# 4.50fF
C45 gnd a_1251_110# 5.70fF
C46 vdd b4 3.60fF
C47 vdd a2 3.60fF
C48 s4 Gnd 49.44fF
C49 a_3066_n134# Gnd 84.66fF
C50 a_3206_n36# Gnd 77.63fF
C51 a_2722_n136# Gnd 84.66fF
C52 s3 Gnd 49.44fF
C53 a_3066_0# Gnd 77.73fF
C54 a_2862_n38# Gnd 77.63fF
C55 a_2083_n136# Gnd 84.66fF
C56 a_3402_44# Gnd 91.16fF
C57 cout Gnd 66.73fF
C58 a_2722_n2# Gnd 77.73fF
C59 a_2223_n38# Gnd 77.63fF
C60 a_1739_n138# Gnd 84.66fF
C61 s2 Gnd 49.12fF
C62 a_2083_n2# Gnd 77.73fF
C63 a_1879_n40# Gnd 77.63fF
C64 a_1061_n138# Gnd 84.66fF
C65 a_2419_42# Gnd 91.16fF
C66 a_3256_114# Gnd 103.86fF
C67 a_3066_154# Gnd 98.68fF
C68 a_2722_152# Gnd 98.68fF
C69 a_2912_112# Gnd 192.16fF
C70 a_2870_n138# Gnd 158.51fF
C71 b4 Gnd 99.91fF
C72 a4 Gnd 99.60fF
C73 a_1739_n4# Gnd 77.73fF
C74 a_1201_n40# Gnd 77.63fF
C75 a_717_n140# Gnd 84.66fF
C76 s1 Gnd 49.12fF
C77 a_1061_n4# Gnd 77.73fF
C78 a_857_n42# Gnd 77.63fF
C79 a_78_n140# Gnd 84.66fF
C80 a_1397_40# Gnd 91.16fF
C81 a_2273_112# Gnd 103.86fF
C82 a_2083_152# Gnd 98.68fF
C83 a_1739_150# Gnd 98.68fF
C84 a_1929_110# Gnd 192.16fF
C85 a_1887_n140# Gnd 158.51fF
C86 b3 Gnd 100.54fF
C87 a3 Gnd 99.60fF
C88 a_717_n6# Gnd 77.73fF
C89 a_218_n42# Gnd 77.63fF
C90 a_n266_n142# Gnd 84.66fF
C91 a_78_n6# Gnd 77.73fF
C92 a_n126_n44# Gnd 77.63fF
C93 a_414_38# Gnd 91.16fF
C94 a_1251_110# Gnd 103.86fF
C95 a_1061_150# Gnd 98.68fF
C96 a_717_148# Gnd 98.68fF
C97 a_907_108# Gnd 192.16fF
C98 a_1575_46# Gnd 381.20fF
C99 a_865_n142# Gnd 158.51fF
C100 b2 Gnd 99.28fF
C101 a2 Gnd 99.28fF
C102 a_n266_n8# Gnd 77.73fF
C103 gnd Gnd 4899.14fF
C104 a_268_108# Gnd 103.86fF
C105 a_78_148# Gnd 98.68fF
C106 a_n266_146# Gnd 98.68fF
C107 vdd Gnd 5079.42fF
C108 a_n76_106# Gnd 192.16fF
C109 cin Gnd 98.65fF
C110 a_n118_n144# Gnd 158.51fF
C111 b1 Gnd 99.28fF
C112 a1 Gnd 99.60fF
C113 a_592_44# Gnd 381.52fF
C114 a_2597_48# Gnd 381.52fF
