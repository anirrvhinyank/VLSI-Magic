magic
tech scmos
timestamp 1635335426
<< nwell >>
rect -9 -1 37 11
<< polysilicon >>
rect -2 9 0 11
rect 8 9 10 11
rect 27 9 29 11
rect -2 -4 0 1
rect -1 -8 0 -4
rect -2 -18 0 -8
rect 8 -10 10 1
rect 27 -3 29 1
rect 20 -7 29 -3
rect 9 -14 10 -10
rect 8 -18 10 -14
rect 27 -18 29 -7
rect -2 -28 0 -26
rect 8 -28 10 -26
rect 27 -28 29 -26
<< ndiffusion >>
rect -7 -20 -2 -18
rect -3 -24 -2 -20
rect -7 -26 -2 -24
rect 0 -26 8 -18
rect 10 -20 17 -18
rect 10 -24 12 -20
rect 16 -24 17 -20
rect 10 -26 17 -24
rect 21 -20 27 -18
rect 25 -24 27 -20
rect 21 -26 27 -24
rect 29 -20 35 -18
rect 29 -24 31 -20
rect 29 -26 35 -24
<< pdiffusion >>
rect -7 7 -2 9
rect -3 3 -2 7
rect -7 1 -2 3
rect 0 7 8 9
rect 0 3 2 7
rect 6 3 8 7
rect 0 1 8 3
rect 10 7 17 9
rect 10 3 12 7
rect 16 3 17 7
rect 10 1 17 3
rect 21 7 27 9
rect 25 3 27 7
rect 21 1 27 3
rect 29 7 35 9
rect 29 3 31 7
rect 29 1 35 3
<< metal1 >>
rect -7 13 2 17
rect 6 13 12 17
rect 16 13 21 17
rect -7 7 -3 13
rect 12 7 16 13
rect 21 7 25 13
rect 2 -3 6 3
rect 31 -3 35 3
rect -6 -8 -5 -4
rect 2 -7 16 -3
rect 31 -7 38 -3
rect 4 -14 5 -10
rect 12 -20 16 -7
rect 31 -20 35 -7
rect -7 -30 -3 -24
rect 21 -30 25 -24
rect -7 -34 2 -30
rect 6 -34 11 -30
rect 15 -34 21 -30
<< ntransistor >>
rect -2 -26 0 -18
rect 8 -26 10 -18
rect 27 -26 29 -18
<< ptransistor >>
rect -2 1 0 9
rect 8 1 10 9
rect 27 1 29 9
<< polycontact >>
rect -5 -8 -1 -4
rect 16 -7 20 -3
rect 5 -14 9 -10
<< ndcontact >>
rect -7 -24 -3 -20
rect 12 -24 16 -20
rect 21 -24 25 -20
rect 31 -24 35 -20
<< pdcontact >>
rect -7 3 -3 7
rect 2 3 6 7
rect 12 3 16 7
rect 21 3 25 7
rect 31 3 35 7
<< psubstratepcontact >>
rect -7 -34 -3 -30
rect 2 -34 6 -30
rect 11 -34 15 -30
rect 21 -34 25 -30
<< nsubstratencontact >>
rect -7 13 -3 17
rect 2 13 6 17
rect 12 13 16 17
rect 21 13 25 17
<< labels >>
rlabel metal1 -2 15 -2 15 5 vdd
rlabel metal1 -2 -32 -2 -32 1 vss
rlabel polycontact -3 -6 -3 -6 1 a
rlabel metal1 34 -5 34 -5 7 out
rlabel polycontact 7 -12 7 -12 1 b
<< end >>
