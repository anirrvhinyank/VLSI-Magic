magic
tech scmos
timestamp 1636294044
<< polysilicon >>
rect -807 700 -210 704
rect -214 698 -210 700
rect -480 651 117 655
rect -875 405 -544 409
rect -875 326 -871 405
rect -807 326 -803 383
rect -685 318 -681 339
rect -548 326 -544 405
rect -480 326 -476 651
rect -282 596 49 600
rect -282 517 -278 596
rect -214 517 -210 571
rect -92 509 -88 530
rect 45 517 49 596
rect 113 517 117 651
rect -282 473 -278 497
rect -214 473 -210 497
rect 235 509 239 519
rect -92 483 -88 489
rect 45 473 49 497
rect 113 473 117 497
rect 235 483 239 489
rect -92 467 -88 473
rect -282 458 -278 463
rect -214 405 -210 463
rect 235 467 239 473
rect 45 458 49 463
rect 113 458 117 463
rect -92 450 -88 457
rect 235 452 239 457
rect -202 351 -148 361
rect -875 282 -871 306
rect -807 282 -803 306
rect -358 318 -354 328
rect -685 292 -681 298
rect -548 282 -544 306
rect -480 282 -476 306
rect -358 292 -354 298
rect -685 276 -681 282
rect -875 267 -871 272
rect -807 267 -803 272
rect -358 276 -354 282
rect -548 267 -544 272
rect -480 267 -476 272
rect -685 259 -681 266
rect -358 261 -354 266
rect -270 166 -266 244
rect -202 166 -198 351
rect 628 295 1129 299
rect 74 168 78 188
rect 142 168 146 228
rect 410 210 414 212
rect 412 200 414 210
rect -80 158 -76 164
rect -270 122 -266 146
rect -202 122 -198 146
rect 264 160 268 166
rect -80 132 -76 138
rect 74 124 78 148
rect 142 124 146 148
rect 264 134 268 140
rect -80 116 -76 122
rect -270 12 -266 112
rect -202 12 -198 112
rect 264 118 268 124
rect -80 100 -76 106
rect -130 8 -126 28
rect 74 14 78 114
rect 142 14 146 114
rect 264 102 268 108
rect 410 92 414 200
rect 628 138 632 295
rect 713 168 717 267
rect 781 168 785 266
rect 1057 170 1061 190
rect 1125 170 1129 295
rect 1393 212 1397 214
rect 1395 202 1397 212
rect 903 160 907 166
rect 713 124 717 148
rect 781 124 785 148
rect 1247 162 1251 168
rect 903 134 907 140
rect 1057 126 1061 150
rect 1125 126 1129 150
rect 1247 136 1251 142
rect 903 118 907 124
rect 478 92 482 112
rect 588 96 592 102
rect 410 48 414 72
rect 478 48 482 72
rect 588 70 592 76
rect 588 54 592 60
rect 588 38 592 44
rect -270 -32 -266 -8
rect -202 -32 -198 -8
rect 214 10 218 30
rect 410 18 414 38
rect 478 16 482 38
rect -130 -18 -126 -12
rect -54 -18 -50 -6
rect -130 -34 -126 -28
rect -270 -88 -266 -42
rect -202 -88 -198 -42
rect -130 -50 -126 -44
rect -122 -90 -118 -70
rect -54 -90 -50 -28
rect 74 -30 78 -6
rect 142 -30 146 -6
rect 713 14 717 114
rect 781 14 785 114
rect 1247 120 1251 126
rect 903 102 907 108
rect 478 4 482 6
rect 214 -16 218 -10
rect 290 -16 294 -4
rect 853 10 857 30
rect 1057 16 1061 116
rect 1125 16 1129 116
rect 1247 104 1251 110
rect 1393 94 1397 202
rect 1611 140 1615 155
rect 1461 94 1465 114
rect 1571 98 1575 104
rect 1393 50 1397 74
rect 1461 50 1465 74
rect 1571 72 1575 78
rect 1571 56 1575 62
rect 1571 40 1575 46
rect 214 -32 218 -26
rect 74 -86 78 -40
rect 142 -86 146 -40
rect 214 -48 218 -42
rect -270 -132 -266 -108
rect -202 -132 -198 -108
rect 222 -88 226 -68
rect 290 -88 294 -26
rect 713 -30 717 -6
rect 781 -30 785 -6
rect 1197 12 1201 32
rect 1393 20 1397 40
rect 1461 18 1465 40
rect 853 -16 857 -10
rect 929 -16 933 -4
rect 853 -32 857 -26
rect 713 -86 717 -40
rect 781 -86 785 -40
rect 853 -48 857 -42
rect -122 -114 -118 -110
rect -122 -134 -118 -124
rect -54 -134 -50 -110
rect 74 -118 78 -106
rect -16 -122 78 -118
rect 74 -130 78 -122
rect 142 -130 146 -106
rect 861 -88 865 -68
rect 929 -88 933 -26
rect 1057 -28 1061 -4
rect 1125 -28 1129 -4
rect 1461 6 1465 8
rect 1197 -14 1201 -8
rect 1273 -14 1277 -2
rect 1197 -30 1201 -24
rect 1057 -84 1061 -38
rect 1125 -84 1129 -38
rect 1197 -46 1201 -40
rect 222 -112 226 -108
rect -270 -162 -266 -142
rect -202 -162 -198 -142
rect 222 -132 226 -122
rect 290 -132 294 -108
rect 328 -120 342 -116
rect 713 -130 717 -106
rect 781 -130 785 -106
rect 1205 -86 1209 -66
rect 1273 -86 1277 -24
rect 861 -112 865 -108
rect -122 -164 -118 -144
rect -54 -164 -50 -144
rect 74 -160 78 -140
rect 142 -160 146 -140
rect 861 -132 865 -122
rect 929 -132 933 -108
rect 1057 -116 1061 -104
rect 967 -120 1061 -116
rect 1057 -128 1061 -120
rect 1125 -128 1129 -104
rect 1205 -110 1209 -106
rect 222 -162 226 -142
rect 290 -162 294 -142
rect 713 -160 717 -140
rect 781 -160 785 -140
rect 1205 -130 1209 -120
rect 1273 -130 1277 -106
rect 1311 -118 1325 -114
rect 861 -162 865 -142
rect 929 -162 933 -142
rect 1057 -158 1061 -138
rect 1125 -158 1129 -138
rect 1205 -160 1209 -140
rect 1273 -160 1277 -140
<< ndiffusion >>
rect -300 463 -298 473
rect -288 463 -282 473
rect -278 463 -214 473
rect -210 463 -206 473
rect -196 463 -194 473
rect -114 457 -112 467
rect -102 457 -92 467
rect -88 457 -78 467
rect -68 457 -66 467
rect 27 463 29 473
rect 39 463 45 473
rect 49 463 113 473
rect 117 463 121 473
rect 131 463 133 473
rect 213 457 215 467
rect 225 457 235 467
rect 239 457 249 467
rect 259 457 261 467
rect -893 272 -891 282
rect -881 272 -875 282
rect -871 272 -807 282
rect -803 272 -799 282
rect -789 272 -787 282
rect -707 266 -705 276
rect -695 266 -685 276
rect -681 266 -671 276
rect -661 266 -659 276
rect -566 272 -564 282
rect -554 272 -548 282
rect -544 272 -480 282
rect -476 272 -472 282
rect -462 272 -460 282
rect -380 266 -378 276
rect -368 266 -358 276
rect -354 266 -344 276
rect -334 266 -332 276
rect -288 112 -286 122
rect -276 112 -270 122
rect -266 112 -202 122
rect -198 112 -194 122
rect -184 112 -182 122
rect -102 106 -100 116
rect -90 106 -80 116
rect -76 106 -66 116
rect -56 106 -54 116
rect 56 114 58 124
rect 68 114 74 124
rect 78 114 142 124
rect 146 114 150 124
rect 160 114 162 124
rect 242 108 244 118
rect 254 108 264 118
rect 268 108 278 118
rect 288 108 290 118
rect 695 114 697 124
rect 707 114 713 124
rect 717 114 781 124
rect 785 114 789 124
rect 799 114 801 124
rect 392 38 394 48
rect 404 38 410 48
rect 414 38 436 48
rect 446 38 478 48
rect 482 38 486 48
rect 496 38 498 48
rect 566 44 568 54
rect 578 44 588 54
rect 592 44 602 54
rect 612 44 614 54
rect -288 -42 -286 -32
rect -276 -42 -270 -32
rect -266 -42 -202 -32
rect -198 -42 -194 -32
rect -184 -42 -182 -32
rect -152 -44 -150 -34
rect -140 -44 -130 -34
rect -126 -44 -116 -34
rect -106 -44 -104 -34
rect 881 108 883 118
rect 893 108 903 118
rect 907 108 917 118
rect 927 108 929 118
rect 1039 116 1041 126
rect 1051 116 1057 126
rect 1061 116 1125 126
rect 1129 116 1133 126
rect 1143 116 1145 126
rect 1225 110 1227 120
rect 1237 110 1247 120
rect 1251 110 1261 120
rect 1271 110 1273 120
rect 1375 40 1377 50
rect 1387 40 1393 50
rect 1397 40 1419 50
rect 1429 40 1461 50
rect 1465 40 1469 50
rect 1479 40 1481 50
rect 1549 46 1551 56
rect 1561 46 1571 56
rect 1575 46 1585 56
rect 1595 46 1597 56
rect 56 -40 58 -30
rect 68 -40 74 -30
rect 78 -40 142 -30
rect 146 -40 150 -30
rect 160 -40 162 -30
rect 192 -42 194 -32
rect 204 -42 214 -32
rect 218 -42 228 -32
rect 238 -42 240 -32
rect 695 -40 697 -30
rect 707 -40 713 -30
rect 717 -40 781 -30
rect 785 -40 789 -30
rect 799 -40 801 -30
rect 831 -42 833 -32
rect 843 -42 853 -32
rect 857 -42 867 -32
rect 877 -42 879 -32
rect -288 -142 -286 -132
rect -276 -142 -270 -132
rect -266 -142 -244 -132
rect -234 -142 -202 -132
rect -198 -142 -194 -132
rect -184 -142 -182 -132
rect 1039 -38 1041 -28
rect 1051 -38 1057 -28
rect 1061 -38 1125 -28
rect 1129 -38 1133 -28
rect 1143 -38 1145 -28
rect 1175 -40 1177 -30
rect 1187 -40 1197 -30
rect 1201 -40 1211 -30
rect 1221 -40 1223 -30
rect -140 -144 -138 -134
rect -128 -144 -122 -134
rect -118 -144 -96 -134
rect -86 -144 -54 -134
rect -50 -144 -46 -134
rect -36 -144 -34 -134
rect 56 -140 58 -130
rect 68 -140 74 -130
rect 78 -140 100 -130
rect 110 -140 142 -130
rect 146 -140 150 -130
rect 160 -140 162 -130
rect 204 -142 206 -132
rect 216 -142 222 -132
rect 226 -142 248 -132
rect 258 -142 290 -132
rect 294 -142 298 -132
rect 308 -142 310 -132
rect 695 -140 697 -130
rect 707 -140 713 -130
rect 717 -140 739 -130
rect 749 -140 781 -130
rect 785 -140 789 -130
rect 799 -140 801 -130
rect 843 -142 845 -132
rect 855 -142 861 -132
rect 865 -142 887 -132
rect 897 -142 929 -132
rect 933 -142 937 -132
rect 947 -142 949 -132
rect 1039 -138 1041 -128
rect 1051 -138 1057 -128
rect 1061 -138 1083 -128
rect 1093 -138 1125 -128
rect 1129 -138 1133 -128
rect 1143 -138 1145 -128
rect 1187 -140 1189 -130
rect 1199 -140 1205 -130
rect 1209 -140 1231 -130
rect 1241 -140 1273 -130
rect 1277 -140 1281 -130
rect 1291 -140 1293 -130
<< pdiffusion >>
rect -893 320 -875 326
rect -893 310 -891 320
rect -881 310 -875 320
rect -893 306 -875 310
rect -871 320 -807 326
rect -871 310 -849 320
rect -839 310 -807 320
rect -871 306 -807 310
rect -803 320 -787 326
rect -803 310 -799 320
rect -789 310 -787 320
rect -300 511 -282 517
rect -300 501 -298 511
rect -288 501 -282 511
rect -300 497 -282 501
rect -278 511 -214 517
rect -278 501 -256 511
rect -246 501 -214 511
rect -278 497 -214 501
rect -210 511 -194 517
rect -210 501 -206 511
rect -196 501 -194 511
rect 27 511 45 517
rect -210 497 -194 501
rect -114 505 -92 509
rect -114 495 -112 505
rect -102 495 -92 505
rect -114 489 -92 495
rect -88 505 -66 509
rect -88 495 -78 505
rect -68 495 -66 505
rect 27 501 29 511
rect 39 501 45 511
rect 27 497 45 501
rect 49 511 113 517
rect 49 501 71 511
rect 81 501 113 511
rect 49 497 113 501
rect 117 511 133 517
rect 117 501 121 511
rect 131 501 133 511
rect 117 497 133 501
rect 213 505 235 509
rect -88 489 -66 495
rect 213 495 215 505
rect 225 495 235 505
rect 213 489 235 495
rect 239 505 261 509
rect 239 495 249 505
rect 259 495 261 505
rect 239 489 261 495
rect -566 320 -548 326
rect -803 306 -787 310
rect -707 314 -685 318
rect -707 304 -705 314
rect -695 304 -685 314
rect -707 298 -685 304
rect -681 314 -659 318
rect -681 304 -671 314
rect -661 304 -659 314
rect -566 310 -564 320
rect -554 310 -548 320
rect -566 306 -548 310
rect -544 320 -480 326
rect -544 310 -522 320
rect -512 310 -480 320
rect -544 306 -480 310
rect -476 320 -460 326
rect -476 310 -472 320
rect -462 310 -460 320
rect -476 306 -460 310
rect -380 314 -358 318
rect -681 298 -659 304
rect -380 304 -378 314
rect -368 304 -358 314
rect -380 298 -358 304
rect -354 314 -332 318
rect -354 304 -344 314
rect -334 304 -332 314
rect -354 298 -332 304
rect -288 160 -270 166
rect -288 150 -286 160
rect -276 150 -270 160
rect -288 146 -270 150
rect -266 160 -202 166
rect -266 150 -244 160
rect -234 150 -202 160
rect -266 146 -202 150
rect -198 160 -182 166
rect -198 150 -194 160
rect -184 150 -182 160
rect 56 162 74 168
rect -198 146 -182 150
rect -102 154 -80 158
rect -102 144 -100 154
rect -90 144 -80 154
rect -102 138 -80 144
rect -76 154 -54 158
rect -76 144 -66 154
rect -56 144 -54 154
rect 56 152 58 162
rect 68 152 74 162
rect 56 148 74 152
rect 78 162 142 168
rect 78 152 100 162
rect 110 152 142 162
rect 78 148 142 152
rect 146 162 162 168
rect 146 152 150 162
rect 160 152 162 162
rect 146 148 162 152
rect 242 156 264 160
rect -76 138 -54 144
rect 242 146 244 156
rect 254 146 264 156
rect 242 140 264 146
rect 268 156 290 160
rect 268 146 278 156
rect 288 146 290 156
rect 268 140 290 146
rect -288 6 -270 12
rect -288 -4 -286 6
rect -276 -4 -270 6
rect -288 -8 -270 -4
rect -266 6 -202 12
rect -266 -4 -244 6
rect -234 -4 -202 6
rect -266 -8 -202 -4
rect -198 6 -182 12
rect 695 162 713 168
rect 695 152 697 162
rect 707 152 713 162
rect 695 148 713 152
rect 717 162 781 168
rect 717 152 739 162
rect 749 152 781 162
rect 717 148 781 152
rect 785 162 801 168
rect 785 152 789 162
rect 799 152 801 162
rect 1039 164 1057 170
rect 785 148 801 152
rect 881 156 903 160
rect 881 146 883 156
rect 893 146 903 156
rect 881 140 903 146
rect 907 156 929 160
rect 907 146 917 156
rect 927 146 929 156
rect 1039 154 1041 164
rect 1051 154 1057 164
rect 1039 150 1057 154
rect 1061 164 1125 170
rect 1061 154 1083 164
rect 1093 154 1125 164
rect 1061 150 1125 154
rect 1129 164 1145 170
rect 1129 154 1133 164
rect 1143 154 1145 164
rect 1129 150 1145 154
rect 1225 158 1247 162
rect 907 140 929 146
rect 1225 148 1227 158
rect 1237 148 1247 158
rect 1225 142 1247 148
rect 1251 158 1273 162
rect 1251 148 1261 158
rect 1271 148 1273 158
rect 1251 142 1273 148
rect 566 92 588 96
rect 392 86 410 92
rect 392 76 394 86
rect 404 76 410 86
rect 392 72 410 76
rect 414 72 478 92
rect 482 86 498 92
rect 482 76 486 86
rect 496 76 498 86
rect 566 82 568 92
rect 578 82 588 92
rect 566 76 588 82
rect 592 92 614 96
rect 592 82 602 92
rect 612 82 614 92
rect 592 76 614 82
rect 482 72 498 76
rect 56 8 74 14
rect -198 -4 -194 6
rect -184 -4 -182 6
rect -198 -8 -182 -4
rect -152 4 -130 8
rect -152 -6 -150 4
rect -140 -6 -130 4
rect -152 -12 -130 -6
rect -126 4 -104 8
rect -126 -6 -116 4
rect -106 -6 -104 4
rect 56 -2 58 8
rect 68 -2 74 8
rect 56 -6 74 -2
rect 78 8 142 14
rect 78 -2 100 8
rect 110 -2 142 8
rect 78 -6 142 -2
rect 146 8 162 14
rect 146 -2 150 8
rect 160 -2 162 8
rect 146 -6 162 -2
rect 192 6 214 10
rect 192 -4 194 6
rect 204 -4 214 6
rect -126 -12 -104 -6
rect -288 -94 -270 -88
rect -288 -104 -286 -94
rect -276 -104 -270 -94
rect -288 -108 -270 -104
rect -266 -108 -202 -88
rect -198 -94 -182 -88
rect 192 -10 214 -4
rect 218 6 240 10
rect 218 -4 228 6
rect 238 -4 240 6
rect 695 8 713 14
rect 695 -2 697 8
rect 707 -2 713 8
rect 218 -10 240 -4
rect 695 -6 713 -2
rect 717 8 781 14
rect 717 -2 739 8
rect 749 -2 781 8
rect 717 -6 781 -2
rect 785 8 801 14
rect 1549 94 1571 98
rect 1375 88 1393 94
rect 1375 78 1377 88
rect 1387 78 1393 88
rect 1375 74 1393 78
rect 1397 74 1461 94
rect 1465 88 1481 94
rect 1465 78 1469 88
rect 1479 78 1481 88
rect 1549 84 1551 94
rect 1561 84 1571 94
rect 1549 78 1571 84
rect 1575 94 1597 98
rect 1575 84 1585 94
rect 1595 84 1597 94
rect 1575 78 1597 84
rect 1465 74 1481 78
rect 1039 10 1057 16
rect 785 -2 789 8
rect 799 -2 801 8
rect 785 -6 801 -2
rect 831 6 853 10
rect 831 -4 833 6
rect 843 -4 853 6
rect -198 -104 -194 -94
rect -184 -104 -182 -94
rect -198 -108 -182 -104
rect -140 -96 -122 -90
rect -140 -106 -138 -96
rect -128 -106 -122 -96
rect -140 -110 -122 -106
rect -118 -110 -54 -90
rect -50 -96 -34 -90
rect -50 -106 -46 -96
rect -36 -106 -34 -96
rect 56 -92 74 -86
rect 56 -102 58 -92
rect 68 -102 74 -92
rect 56 -106 74 -102
rect 78 -106 142 -86
rect 146 -92 162 -86
rect 831 -10 853 -4
rect 857 6 879 10
rect 857 -4 867 6
rect 877 -4 879 6
rect 1039 0 1041 10
rect 1051 0 1057 10
rect 1039 -4 1057 0
rect 1061 10 1125 16
rect 1061 0 1083 10
rect 1093 0 1125 10
rect 1061 -4 1125 0
rect 1129 10 1145 16
rect 1129 0 1133 10
rect 1143 0 1145 10
rect 1129 -4 1145 0
rect 1175 8 1197 12
rect 1175 -2 1177 8
rect 1187 -2 1197 8
rect 857 -10 879 -4
rect 146 -102 150 -92
rect 160 -102 162 -92
rect 146 -106 162 -102
rect 204 -94 222 -88
rect 204 -104 206 -94
rect 216 -104 222 -94
rect -50 -110 -34 -106
rect 204 -108 222 -104
rect 226 -108 290 -88
rect 294 -94 310 -88
rect 294 -104 298 -94
rect 308 -104 310 -94
rect 294 -108 310 -104
rect 695 -92 713 -86
rect 695 -102 697 -92
rect 707 -102 713 -92
rect 695 -106 713 -102
rect 717 -106 781 -86
rect 785 -92 801 -86
rect 1175 -8 1197 -2
rect 1201 8 1223 12
rect 1201 -2 1211 8
rect 1221 -2 1223 8
rect 1201 -8 1223 -2
rect 785 -102 789 -92
rect 799 -102 801 -92
rect 785 -106 801 -102
rect 843 -94 861 -88
rect 843 -104 845 -94
rect 855 -104 861 -94
rect 843 -108 861 -104
rect 865 -108 929 -88
rect 933 -94 949 -88
rect 933 -104 937 -94
rect 947 -104 949 -94
rect 1039 -90 1057 -84
rect 1039 -100 1041 -90
rect 1051 -100 1057 -90
rect 1039 -104 1057 -100
rect 1061 -104 1125 -84
rect 1129 -90 1145 -84
rect 1129 -100 1133 -90
rect 1143 -100 1145 -90
rect 1129 -104 1145 -100
rect 1187 -92 1205 -86
rect 1187 -102 1189 -92
rect 1199 -102 1205 -92
rect 933 -108 949 -104
rect 1187 -106 1205 -102
rect 1209 -106 1273 -86
rect 1277 -92 1293 -86
rect 1277 -102 1281 -92
rect 1291 -102 1293 -92
rect 1277 -106 1293 -102
<< metal1 >>
rect -807 387 -803 696
rect -214 575 -210 694
rect 29 554 167 559
rect -420 553 -405 554
rect -114 553 167 554
rect -420 547 167 553
rect 179 547 225 559
rect -420 542 39 547
rect -420 541 -102 542
rect -420 368 -405 541
rect -298 511 -288 541
rect -206 511 -196 541
rect -112 505 -102 541
rect 29 511 39 542
rect 121 511 131 547
rect -256 491 -246 501
rect 215 505 225 547
rect -256 483 -176 491
rect -78 483 -68 495
rect 71 491 81 501
rect 71 483 151 491
rect 249 483 259 495
rect -256 481 -98 483
rect -206 473 -196 481
rect -186 473 -98 481
rect -78 473 -60 483
rect 71 481 229 483
rect 121 473 131 481
rect 141 473 229 481
rect 249 473 267 483
rect -78 467 -68 473
rect -298 435 -288 463
rect 249 467 259 473
rect -112 436 -102 457
rect 29 436 39 463
rect -112 435 39 436
rect -298 433 39 435
rect 215 433 225 457
rect -298 426 225 433
rect -564 362 -368 368
rect -891 356 -368 362
rect -891 351 -554 356
rect -891 350 -695 351
rect -891 320 -881 350
rect -799 320 -789 350
rect -705 314 -695 350
rect -564 320 -554 351
rect -472 320 -462 356
rect -849 300 -839 310
rect -378 314 -368 356
rect -849 292 -769 300
rect -671 292 -661 304
rect -522 300 -512 310
rect -522 292 -442 300
rect -344 292 -334 304
rect -849 290 -691 292
rect -799 282 -789 290
rect -779 282 -691 290
rect -671 282 -653 292
rect -522 290 -364 292
rect -472 282 -462 290
rect -452 282 -364 290
rect -344 282 -326 292
rect -671 276 -661 282
rect -891 244 -881 272
rect -344 276 -334 282
rect -705 245 -695 266
rect -564 245 -554 272
rect -705 244 -554 245
rect -891 242 -554 244
rect -378 242 -368 266
rect -298 242 -288 426
rect 29 424 225 426
rect -138 351 -91 361
rect -270 248 -266 269
rect 713 271 717 400
rect -891 235 -288 242
rect -891 89 -881 235
rect -564 233 -288 235
rect 336 200 402 210
rect 1319 202 1385 212
rect 959 180 1512 182
rect -24 178 1512 180
rect -298 168 -138 178
rect -125 172 1512 178
rect -125 170 969 172
rect -125 168 -14 170
rect -286 160 -276 168
rect -194 160 -184 168
rect -100 154 -90 168
rect -244 140 -234 150
rect -244 132 -164 140
rect -66 132 -56 144
rect -244 130 -86 132
rect -194 122 -184 130
rect -174 122 -86 130
rect -66 122 -48 132
rect -66 116 -56 122
rect -286 106 -276 112
rect -310 100 -164 106
rect -100 100 -90 106
rect -310 96 -90 100
rect -310 89 -300 96
rect -174 90 -90 96
rect -891 77 -300 89
rect -310 -48 -300 77
rect -24 24 -14 168
rect 58 162 68 170
rect 150 162 160 170
rect 244 156 254 170
rect 100 142 110 152
rect 100 134 180 142
rect 278 134 288 146
rect 100 132 258 134
rect 150 124 160 132
rect 170 124 258 132
rect 278 124 296 134
rect 278 118 288 124
rect 58 108 68 114
rect -286 14 -14 24
rect -286 6 -276 14
rect -194 6 -184 14
rect -150 12 -14 14
rect -150 4 -140 12
rect -244 -14 -234 -4
rect -244 -18 -164 -14
rect -116 -18 -106 -6
rect -244 -24 -136 -18
rect -194 -32 -184 -24
rect -174 -28 -136 -24
rect -116 -28 -60 -18
rect -116 -34 -106 -28
rect -286 -48 -276 -42
rect -150 -48 -140 -44
rect -310 -58 -140 -48
rect -310 -150 -300 -58
rect -24 -76 -14 12
rect -286 -86 -14 -76
rect 34 102 180 108
rect 244 102 254 108
rect 34 98 254 102
rect 34 -46 44 98
rect 170 92 254 98
rect 320 104 330 170
rect 697 162 707 170
rect 789 162 799 170
rect 883 156 893 170
rect 739 142 749 152
rect 739 134 819 142
rect 917 134 927 146
rect 739 132 897 134
rect 394 104 578 106
rect 392 96 578 104
rect 392 94 404 96
rect 320 26 330 94
rect 394 86 404 94
rect 568 92 578 96
rect 486 66 496 76
rect 602 70 612 82
rect 624 70 634 128
rect 789 124 799 132
rect 809 124 897 132
rect 917 124 935 134
rect 917 118 927 124
rect 697 108 707 114
rect 506 66 582 70
rect 436 60 582 66
rect 602 60 634 70
rect 673 102 819 108
rect 883 102 893 108
rect 673 98 893 102
rect 436 56 516 60
rect 436 48 446 56
rect 602 54 612 60
rect 58 16 330 26
rect 58 8 68 16
rect 150 8 160 16
rect 194 14 330 16
rect 194 6 204 14
rect 100 -12 110 -2
rect 100 -16 180 -12
rect 228 -16 238 -4
rect 100 -22 208 -16
rect 150 -30 160 -22
rect 170 -26 208 -22
rect 228 -26 284 -16
rect 228 -32 238 -26
rect 58 -46 68 -40
rect 194 -46 204 -42
rect 34 -56 204 -46
rect -286 -94 -276 -86
rect -194 -114 -184 -104
rect -138 -96 -128 -86
rect -244 -124 -128 -114
rect -46 -116 -36 -106
rect -244 -132 -234 -124
rect -96 -126 -26 -116
rect -96 -134 -86 -126
rect -286 -150 -276 -142
rect -194 -150 -184 -142
rect -138 -150 -128 -144
rect -46 -150 -36 -144
rect 34 -148 44 -56
rect 320 -74 330 14
rect 58 -84 330 -74
rect 394 32 404 38
rect 486 32 496 38
rect 568 32 578 44
rect 394 22 578 32
rect 58 -92 68 -84
rect 150 -112 160 -102
rect 206 -94 216 -84
rect 100 -122 216 -112
rect 298 -114 308 -104
rect 100 -130 110 -122
rect 248 -124 318 -114
rect 248 -132 258 -124
rect 58 -148 68 -140
rect 150 -148 160 -140
rect 206 -148 216 -142
rect 298 -148 308 -142
rect 394 -148 404 22
rect 516 20 578 22
rect 454 6 472 16
rect 673 -46 683 98
rect 809 92 893 98
rect 959 26 969 170
rect 1041 164 1051 172
rect 1133 164 1143 172
rect 1227 158 1237 172
rect 1083 144 1093 154
rect 1083 136 1163 144
rect 1261 136 1271 148
rect 1083 134 1241 136
rect 1133 126 1143 134
rect 1153 126 1241 134
rect 1261 126 1279 136
rect 1261 120 1271 126
rect 1041 110 1051 116
rect 697 16 969 26
rect 697 8 707 16
rect 789 8 799 16
rect 833 14 969 16
rect 833 6 843 14
rect 739 -12 749 -2
rect 739 -16 819 -12
rect 867 -16 877 -4
rect 739 -22 847 -16
rect 789 -30 799 -22
rect 809 -26 847 -22
rect 867 -26 923 -16
rect 867 -32 877 -26
rect 697 -46 707 -40
rect 833 -46 843 -42
rect 673 -56 843 -46
rect 673 -148 683 -56
rect 959 -74 969 14
rect 697 -84 969 -74
rect 1017 104 1163 110
rect 1227 104 1237 110
rect 1017 100 1237 104
rect 1017 -44 1027 100
rect 1153 94 1237 100
rect 1303 106 1313 172
rect 1377 106 1561 108
rect 1375 98 1561 106
rect 1375 96 1387 98
rect 1303 28 1313 96
rect 1377 88 1387 96
rect 1551 94 1561 98
rect 1469 68 1479 78
rect 1585 72 1595 84
rect 1607 72 1617 130
rect 1489 68 1565 72
rect 1419 62 1565 68
rect 1585 62 1617 72
rect 1419 58 1499 62
rect 1419 50 1429 58
rect 1585 56 1595 62
rect 1041 18 1313 28
rect 1041 10 1051 18
rect 1133 10 1143 18
rect 1177 16 1313 18
rect 1177 8 1187 16
rect 1083 -10 1093 0
rect 1083 -14 1163 -10
rect 1211 -14 1221 -2
rect 1083 -20 1191 -14
rect 1133 -28 1143 -20
rect 1153 -24 1191 -20
rect 1211 -24 1267 -14
rect 1211 -30 1221 -24
rect 1041 -44 1051 -38
rect 1177 -44 1187 -40
rect 1017 -54 1187 -44
rect 697 -92 707 -84
rect 789 -112 799 -102
rect 845 -94 855 -84
rect 739 -122 855 -112
rect 937 -114 947 -104
rect 739 -130 749 -122
rect 887 -124 957 -114
rect 887 -132 897 -124
rect 697 -148 707 -140
rect 789 -148 799 -140
rect 845 -148 855 -142
rect 937 -148 947 -142
rect 1017 -146 1027 -54
rect 1303 -72 1313 16
rect 1041 -82 1313 -72
rect 1377 34 1387 40
rect 1469 34 1479 40
rect 1551 34 1561 46
rect 1377 24 1561 34
rect 1041 -90 1051 -82
rect 1133 -110 1143 -100
rect 1189 -92 1199 -82
rect 1083 -120 1199 -110
rect 1281 -112 1291 -102
rect 1083 -128 1093 -120
rect 1231 -122 1301 -112
rect 1231 -130 1241 -122
rect 1041 -146 1051 -138
rect 1133 -146 1143 -138
rect 1189 -146 1199 -140
rect 1281 -146 1291 -140
rect 1377 -146 1387 24
rect 1499 22 1561 24
rect 1437 8 1455 18
rect 1017 -148 1391 -146
rect 34 -150 1391 -148
rect -310 -156 1391 -150
rect -310 -158 1027 -156
rect -310 -160 44 -158
<< metal2 >>
rect -50 473 -30 483
rect -39 361 -30 473
rect -81 351 -30 361
rect 167 409 178 547
rect 283 483 286 518
rect 277 473 286 483
rect 167 320 179 409
rect 717 400 1730 404
rect -138 309 179 320
rect -643 282 -623 292
rect -316 282 -266 292
rect -632 76 -623 282
rect -270 273 -266 282
rect -138 178 -125 309
rect -32 200 326 210
rect 951 202 1309 212
rect -32 132 -22 200
rect 951 134 961 202
rect -38 122 -22 132
rect 945 124 961 134
rect -633 26 -623 76
rect -633 -236 -624 26
rect 296 16 306 124
rect 330 94 382 104
rect 1279 18 1289 126
rect 1313 96 1365 106
rect 296 6 444 16
rect 472 6 482 16
rect 1279 8 1427 18
rect 1455 8 1465 18
rect -632 -249 -624 -236
rect 1712 -249 1730 400
rect -632 -267 1730 -249
rect -632 -268 1704 -267
<< ntransistor >>
rect -282 463 -278 473
rect -214 463 -210 473
rect -92 457 -88 467
rect 45 463 49 473
rect 113 463 117 473
rect 235 457 239 467
rect -875 272 -871 282
rect -807 272 -803 282
rect -685 266 -681 276
rect -548 272 -544 282
rect -480 272 -476 282
rect -358 266 -354 276
rect -270 112 -266 122
rect -202 112 -198 122
rect -80 106 -76 116
rect 74 114 78 124
rect 142 114 146 124
rect 264 108 268 118
rect 713 114 717 124
rect 781 114 785 124
rect 410 38 414 48
rect 478 38 482 48
rect 588 44 592 54
rect -270 -42 -266 -32
rect -202 -42 -198 -32
rect -130 -44 -126 -34
rect 903 108 907 118
rect 1057 116 1061 126
rect 1125 116 1129 126
rect 1247 110 1251 120
rect 1393 40 1397 50
rect 1461 40 1465 50
rect 1571 46 1575 56
rect 74 -40 78 -30
rect 142 -40 146 -30
rect 214 -42 218 -32
rect 713 -40 717 -30
rect 781 -40 785 -30
rect 853 -42 857 -32
rect -270 -142 -266 -132
rect -202 -142 -198 -132
rect 1057 -38 1061 -28
rect 1125 -38 1129 -28
rect 1197 -40 1201 -30
rect -122 -144 -118 -134
rect -54 -144 -50 -134
rect 74 -140 78 -130
rect 142 -140 146 -130
rect 222 -142 226 -132
rect 290 -142 294 -132
rect 713 -140 717 -130
rect 781 -140 785 -130
rect 861 -142 865 -132
rect 929 -142 933 -132
rect 1057 -138 1061 -128
rect 1125 -138 1129 -128
rect 1205 -140 1209 -130
rect 1273 -140 1277 -130
<< ptransistor >>
rect -875 306 -871 326
rect -807 306 -803 326
rect -282 497 -278 517
rect -214 497 -210 517
rect -92 489 -88 509
rect 45 497 49 517
rect 113 497 117 517
rect 235 489 239 509
rect -685 298 -681 318
rect -548 306 -544 326
rect -480 306 -476 326
rect -358 298 -354 318
rect -270 146 -266 166
rect -202 146 -198 166
rect -80 138 -76 158
rect 74 148 78 168
rect 142 148 146 168
rect 264 140 268 160
rect -270 -8 -266 12
rect -202 -8 -198 12
rect 713 148 717 168
rect 781 148 785 168
rect 903 140 907 160
rect 1057 150 1061 170
rect 1125 150 1129 170
rect 1247 142 1251 162
rect 410 72 414 92
rect 478 72 482 92
rect 588 76 592 96
rect -130 -12 -126 8
rect 74 -6 78 14
rect 142 -6 146 14
rect -270 -108 -266 -88
rect -202 -108 -198 -88
rect 214 -10 218 10
rect 713 -6 717 14
rect 781 -6 785 14
rect 1393 74 1397 94
rect 1461 74 1465 94
rect 1571 78 1575 98
rect -122 -110 -118 -90
rect -54 -110 -50 -90
rect 74 -106 78 -86
rect 142 -106 146 -86
rect 853 -10 857 10
rect 1057 -4 1061 16
rect 1125 -4 1129 16
rect 222 -108 226 -88
rect 290 -108 294 -88
rect 713 -106 717 -86
rect 781 -106 785 -86
rect 1197 -8 1201 12
rect 861 -108 865 -88
rect 929 -108 933 -88
rect 1057 -104 1061 -84
rect 1125 -104 1129 -84
rect 1205 -106 1209 -86
rect 1273 -106 1277 -86
<< polycontact >>
rect -807 696 -803 700
rect -214 694 -210 698
rect -807 383 -803 387
rect -214 571 -210 575
rect -98 473 -88 483
rect 229 473 239 483
rect -148 351 -138 361
rect -691 282 -681 292
rect -364 282 -354 292
rect -270 244 -266 248
rect 402 200 412 210
rect -86 122 -76 132
rect 258 124 268 134
rect 713 267 717 271
rect 1385 202 1395 212
rect 624 128 634 138
rect 897 124 907 134
rect 1241 126 1251 136
rect 582 60 592 70
rect -136 -28 -126 -18
rect -60 -28 -50 -18
rect 472 6 482 16
rect 1607 130 1617 140
rect 1565 62 1575 72
rect 208 -26 218 -16
rect 284 -26 294 -16
rect 847 -26 857 -16
rect 923 -26 933 -16
rect -128 -124 -118 -114
rect -26 -126 -16 -116
rect 1455 8 1465 18
rect 1191 -24 1201 -14
rect 1267 -24 1277 -14
rect 216 -122 226 -112
rect 318 -124 328 -114
rect 855 -122 865 -112
rect 957 -124 967 -114
rect 1199 -120 1209 -110
rect 1301 -122 1311 -112
<< ndcontact >>
rect -298 463 -288 473
rect -206 463 -196 473
rect -112 457 -102 467
rect -78 457 -68 467
rect 29 463 39 473
rect 121 463 131 473
rect 215 457 225 467
rect 249 457 259 467
rect -891 272 -881 282
rect -799 272 -789 282
rect -705 266 -695 276
rect -671 266 -661 276
rect -564 272 -554 282
rect -472 272 -462 282
rect -378 266 -368 276
rect -344 266 -334 276
rect -286 112 -276 122
rect -194 112 -184 122
rect -100 106 -90 116
rect -66 106 -56 116
rect 58 114 68 124
rect 150 114 160 124
rect 244 108 254 118
rect 278 108 288 118
rect 697 114 707 124
rect 789 114 799 124
rect 394 38 404 48
rect 436 38 446 48
rect 486 38 496 48
rect 568 44 578 54
rect 602 44 612 54
rect -286 -42 -276 -32
rect -194 -42 -184 -32
rect -150 -44 -140 -34
rect -116 -44 -106 -34
rect 883 108 893 118
rect 917 108 927 118
rect 1041 116 1051 126
rect 1133 116 1143 126
rect 1227 110 1237 120
rect 1261 110 1271 120
rect 1377 40 1387 50
rect 1419 40 1429 50
rect 1469 40 1479 50
rect 1551 46 1561 56
rect 1585 46 1595 56
rect 58 -40 68 -30
rect 150 -40 160 -30
rect 194 -42 204 -32
rect 228 -42 238 -32
rect 697 -40 707 -30
rect 789 -40 799 -30
rect 833 -42 843 -32
rect 867 -42 877 -32
rect -286 -142 -276 -132
rect -244 -142 -234 -132
rect -194 -142 -184 -132
rect 1041 -38 1051 -28
rect 1133 -38 1143 -28
rect 1177 -40 1187 -30
rect 1211 -40 1221 -30
rect -138 -144 -128 -134
rect -96 -144 -86 -134
rect -46 -144 -36 -134
rect 58 -140 68 -130
rect 100 -140 110 -130
rect 150 -140 160 -130
rect 206 -142 216 -132
rect 248 -142 258 -132
rect 298 -142 308 -132
rect 697 -140 707 -130
rect 739 -140 749 -130
rect 789 -140 799 -130
rect 845 -142 855 -132
rect 887 -142 897 -132
rect 937 -142 947 -132
rect 1041 -138 1051 -128
rect 1083 -138 1093 -128
rect 1133 -138 1143 -128
rect 1189 -140 1199 -130
rect 1231 -140 1241 -130
rect 1281 -140 1291 -130
<< pdcontact >>
rect -891 310 -881 320
rect -849 310 -839 320
rect -799 310 -789 320
rect -298 501 -288 511
rect -256 501 -246 511
rect -206 501 -196 511
rect -112 495 -102 505
rect -78 495 -68 505
rect 29 501 39 511
rect 71 501 81 511
rect 121 501 131 511
rect 215 495 225 505
rect 249 495 259 505
rect -705 304 -695 314
rect -671 304 -661 314
rect -564 310 -554 320
rect -522 310 -512 320
rect -472 310 -462 320
rect -378 304 -368 314
rect -344 304 -334 314
rect -286 150 -276 160
rect -244 150 -234 160
rect -194 150 -184 160
rect -100 144 -90 154
rect -66 144 -56 154
rect 58 152 68 162
rect 100 152 110 162
rect 150 152 160 162
rect 244 146 254 156
rect 278 146 288 156
rect -286 -4 -276 6
rect -244 -4 -234 6
rect 697 152 707 162
rect 739 152 749 162
rect 789 152 799 162
rect 883 146 893 156
rect 917 146 927 156
rect 1041 154 1051 164
rect 1083 154 1093 164
rect 1133 154 1143 164
rect 1227 148 1237 158
rect 1261 148 1271 158
rect 394 76 404 86
rect 486 76 496 86
rect 568 82 578 92
rect 602 82 612 92
rect -194 -4 -184 6
rect -150 -6 -140 4
rect -116 -6 -106 4
rect 58 -2 68 8
rect 100 -2 110 8
rect 150 -2 160 8
rect 194 -4 204 6
rect -286 -104 -276 -94
rect 228 -4 238 6
rect 697 -2 707 8
rect 739 -2 749 8
rect 1377 78 1387 88
rect 1469 78 1479 88
rect 1551 84 1561 94
rect 1585 84 1595 94
rect 789 -2 799 8
rect 833 -4 843 6
rect -194 -104 -184 -94
rect -138 -106 -128 -96
rect -46 -106 -36 -96
rect 58 -102 68 -92
rect 867 -4 877 6
rect 1041 0 1051 10
rect 1083 0 1093 10
rect 1133 0 1143 10
rect 1177 -2 1187 8
rect 150 -102 160 -92
rect 206 -104 216 -94
rect 298 -104 308 -94
rect 697 -102 707 -92
rect 1211 -2 1221 8
rect 789 -102 799 -92
rect 845 -104 855 -94
rect 937 -104 947 -94
rect 1041 -100 1051 -90
rect 1133 -100 1143 -90
rect 1189 -102 1199 -92
rect 1281 -102 1291 -92
<< m2contact >>
rect 167 547 179 559
rect -60 473 -50 483
rect 267 473 277 483
rect -653 282 -643 292
rect -326 282 -316 292
rect 713 400 717 404
rect -91 351 -81 361
rect -270 269 -266 273
rect 326 200 336 210
rect 1309 202 1319 212
rect -138 168 -125 178
rect -48 122 -38 132
rect 296 124 306 134
rect 320 94 330 104
rect 382 94 392 104
rect 935 124 945 134
rect 444 6 454 16
rect 1279 126 1289 136
rect 1303 96 1313 106
rect 1365 96 1375 106
rect 1427 8 1437 18
<< labels >>
rlabel metal1 -305 101 -305 101 3 gnd
rlabel metal1 -291 173 -291 173 1 vdd
rlabel polysilicon 144 224 144 224 5 cin
rlabel polysilicon 715 226 715 226 1 a2
rlabel polysilicon 783 227 783 227 1 b2
rlabel polysilicon -267 223 -267 223 1 a1
rlabel polysilicon -200 222 -200 222 1 b1
rlabel metal2 285 506 285 506 1 P0
rlabel polysilicon -873 377 -873 377 1 B1
rlabel polysilicon -805 377 -805 377 1 A1
rlabel polysilicon -478 395 -478 395 1 A0
rlabel polysilicon -280 567 -280 567 1 B0
rlabel polysilicon 338 -118 338 -118 1 P1
rlabel polysilicon 1322 -116 1322 -116 1 P2
rlabel polysilicon 1613 150 1613 150 1 P3
<< end >>
