magic
tech scmos
timestamp 1635503028
<< nwell >>
rect -1 23 25 35
rect 34 16 50 28
rect -1 -45 25 -33
rect 36 -52 51 -40
rect -1 -108 25 -96
rect 36 -108 63 -96
<< polysilicon >>
rect 6 33 8 47
rect 16 33 18 47
rect 41 26 43 35
rect 6 8 8 25
rect 16 8 18 25
rect 41 15 43 18
rect 39 11 43 15
rect 41 8 43 11
rect 6 -35 8 0
rect 16 -35 18 0
rect 41 -2 43 0
rect 42 -42 44 -33
rect 6 -60 8 -43
rect 16 -60 18 -43
rect 42 -53 44 -50
rect 54 -53 56 -49
rect 40 -57 44 -53
rect 42 -60 44 -57
rect 6 -98 8 -68
rect 16 -98 18 -68
rect 42 -70 44 -68
rect 43 -98 45 -94
rect 54 -98 56 -57
rect 6 -123 8 -106
rect 16 -123 18 -106
rect 43 -114 45 -106
rect 40 -118 45 -114
rect 43 -123 45 -118
rect 54 -123 56 -106
rect 69 -118 76 -114
rect 6 -134 8 -131
rect 16 -134 18 -131
rect 43 -133 45 -131
rect 54 -133 56 -131
<< ndiffusion >>
rect 1 6 6 8
rect 5 2 6 6
rect 1 0 6 2
rect 8 0 16 8
rect 18 6 23 8
rect 18 2 19 6
rect 18 0 23 2
rect 36 6 41 8
rect 40 2 41 6
rect 36 0 41 2
rect 43 6 48 8
rect 43 2 44 6
rect 43 0 48 2
rect 1 -62 6 -60
rect 5 -66 6 -62
rect 1 -68 6 -66
rect 8 -68 16 -60
rect 18 -62 23 -60
rect 18 -66 19 -62
rect 18 -68 23 -66
rect 37 -62 42 -60
rect 41 -66 42 -62
rect 37 -68 42 -66
rect 44 -62 49 -60
rect 44 -66 45 -62
rect 44 -68 49 -66
rect 1 -125 6 -123
rect 5 -129 6 -125
rect 1 -131 6 -129
rect 8 -125 16 -123
rect 8 -129 10 -125
rect 14 -129 16 -125
rect 8 -131 16 -129
rect 18 -125 23 -123
rect 18 -129 19 -125
rect 18 -131 23 -129
rect 38 -125 43 -123
rect 42 -129 43 -125
rect 38 -131 43 -129
rect 45 -125 54 -123
rect 45 -129 47 -125
rect 51 -129 54 -125
rect 45 -131 54 -129
rect 56 -125 61 -123
rect 56 -129 57 -125
rect 56 -131 61 -129
<< pdiffusion >>
rect 1 31 6 33
rect 5 27 6 31
rect 1 25 6 27
rect 8 31 16 33
rect 8 27 10 31
rect 14 27 16 31
rect 8 25 16 27
rect 18 31 23 33
rect 18 27 19 31
rect 18 25 23 27
rect 36 24 41 26
rect 40 20 41 24
rect 36 18 41 20
rect 43 24 48 26
rect 43 20 44 24
rect 43 18 48 20
rect 1 -37 6 -35
rect 5 -41 6 -37
rect 1 -43 6 -41
rect 8 -37 16 -35
rect 8 -41 10 -37
rect 14 -41 16 -37
rect 8 -43 16 -41
rect 18 -37 23 -35
rect 18 -41 19 -37
rect 18 -43 23 -41
rect 37 -44 42 -42
rect 41 -48 42 -44
rect 37 -50 42 -48
rect 44 -44 49 -42
rect 44 -48 45 -44
rect 44 -50 49 -48
rect 1 -100 6 -98
rect 5 -104 6 -100
rect 1 -106 6 -104
rect 8 -106 16 -98
rect 18 -100 23 -98
rect 18 -104 19 -100
rect 18 -106 23 -104
rect 38 -100 43 -98
rect 42 -104 43 -100
rect 38 -106 43 -104
rect 45 -106 54 -98
rect 56 -100 61 -98
rect 56 -104 57 -100
rect 56 -106 61 -104
<< metal1 >>
rect -10 36 79 40
rect 1 31 5 36
rect 19 31 23 36
rect 10 15 14 27
rect 36 24 40 36
rect 44 15 48 20
rect 10 11 35 15
rect 44 11 52 15
rect 19 6 23 11
rect 44 6 48 11
rect 1 -11 5 2
rect 36 -11 40 2
rect -8 -15 40 -11
rect -8 -75 -4 -15
rect 75 -23 79 36
rect 1 -27 79 -23
rect 1 -37 5 -27
rect 19 -37 23 -27
rect 10 -53 14 -41
rect 37 -44 41 -27
rect 45 -53 49 -48
rect 10 -57 36 -53
rect 45 -57 52 -53
rect 19 -62 23 -57
rect 45 -62 49 -57
rect 1 -75 5 -66
rect 37 -75 41 -66
rect -8 -79 41 -75
rect -8 -137 -4 -79
rect 75 -88 79 -27
rect 1 -92 79 -88
rect 1 -100 5 -92
rect 38 -100 42 -92
rect 19 -114 23 -104
rect 57 -114 61 -104
rect 10 -118 36 -114
rect 47 -118 65 -114
rect 10 -125 14 -118
rect 47 -125 51 -118
rect 1 -137 5 -129
rect 19 -137 23 -129
rect 38 -137 42 -129
rect 57 -137 61 -129
rect -8 -141 61 -137
<< ntransistor >>
rect 6 0 8 8
rect 16 0 18 8
rect 41 0 43 8
rect 6 -68 8 -60
rect 16 -68 18 -60
rect 42 -68 44 -60
rect 6 -131 8 -123
rect 16 -131 18 -123
rect 43 -131 45 -123
rect 54 -131 56 -123
<< ptransistor >>
rect 6 25 8 33
rect 16 25 18 33
rect 41 18 43 26
rect 6 -43 8 -35
rect 16 -43 18 -35
rect 42 -50 44 -42
rect 6 -106 8 -98
rect 16 -106 18 -98
rect 43 -106 45 -98
rect 54 -106 56 -98
<< polycontact >>
rect 35 11 39 15
rect 36 -57 40 -53
rect 52 -57 56 -53
rect 36 -118 40 -114
rect 65 -118 69 -114
<< ndcontact >>
rect 1 2 5 6
rect 19 2 23 6
rect 36 2 40 6
rect 44 2 48 6
rect 1 -66 5 -62
rect 19 -66 23 -62
rect 37 -66 41 -62
rect 45 -66 49 -62
rect 1 -129 5 -125
rect 10 -129 14 -125
rect 19 -129 23 -125
rect 38 -129 42 -125
rect 47 -129 51 -125
rect 57 -129 61 -125
<< pdcontact >>
rect 1 27 5 31
rect 10 27 14 31
rect 19 27 23 31
rect 36 20 40 24
rect 44 20 48 24
rect 1 -41 5 -37
rect 10 -41 14 -37
rect 19 -41 23 -37
rect 37 -48 41 -44
rect 45 -48 49 -44
rect 1 -104 5 -100
rect 19 -104 23 -100
rect 38 -104 42 -100
rect 57 -104 61 -100
<< labels >>
rlabel metal1 -8 38 -8 38 3 vdd
rlabel polysilicon 7 45 7 45 5 a
rlabel polysilicon 17 45 17 45 5 b
rlabel metal1 35 -139 35 -139 1 gnd
rlabel polysilicon 72 -116 72 -116 1 sum
rlabel metal1 48 13 48 13 1 carryout
<< end >>
