* SPICE3 file created from 2x4decode.ext - technology: scmos

.option scale=1u

M1000 vdd a0 a_74_n107# w_62_n109# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 a_74_n107# a0 a_74_n129# Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_88_n42# a0' a_74_n42# w_62_n44# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vdd a0 a_74_n243# w_62_n245# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_74_n171# a1 vdd w_62_n173# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_74_n243# a0 a_74_n265# Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_74_n42# a0' a_74_n64# Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_74_n193# a1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a1' a1 vdd w_n21_1# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a0' a0 vdd w_27_2# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_74_n107# a1' vdd w_62_n109# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_74_n129# a1' gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 a_74_n243# a1 vdd w_62_n245# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 a_74_n265# a1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 a0' a0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 d2 a_74_n171# vdd w_62_n173# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 d2 a_74_n171# gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 d0 a_74_n42# vdd w_62_n44# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 a1' a1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 d0 a_74_n42# gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 a_74_n42# a1' vdd w_62_n44# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 a_74_n64# a1' gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 d1 a_74_n107# vdd w_62_n109# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 d1 a_74_n107# gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 d3 a_74_n243# vdd w_62_n245# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 vdd a_86_n195# a_74_n171# w_62_n173# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 d3 a_74_n243# gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 a_74_n171# a_86_n195# a_74_n193# Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 d3 Gnd 3.76fF
C1 a_74_n243# Gnd 14.11fF
C2 d2 Gnd 3.76fF
C3 a_74_n171# Gnd 14.11fF
C4 a_86_n195# Gnd 38.96fF
C5 d1 Gnd 3.76fF
C6 a_74_n107# Gnd 14.11fF
C7 d0 Gnd 3.76fF
C8 a_74_n42# Gnd 14.59fF
C9 gnd Gnd 169.00fF
C10 a0' Gnd 46.08fF
C11 a1' Gnd 56.46fF
C12 vdd Gnd 194.39fF
C13 a0 Gnd 66.03fF
C14 a1 Gnd 105.59fF
