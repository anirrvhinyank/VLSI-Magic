magic
tech scmos
timestamp 1636139167
<< polysilicon >>
rect 2633 299 3134 303
rect 628 295 1129 299
rect -270 166 -266 229
rect -202 166 -198 228
rect 74 168 78 188
rect 142 168 146 228
rect 410 210 414 212
rect 412 200 414 210
rect -80 158 -76 164
rect -270 122 -266 146
rect -202 122 -198 146
rect 264 160 268 166
rect -80 132 -76 138
rect 74 124 78 148
rect 142 124 146 148
rect 264 134 268 140
rect -80 116 -76 122
rect -270 12 -266 112
rect -202 12 -198 112
rect 264 118 268 124
rect -80 100 -76 106
rect -130 8 -126 28
rect 74 14 78 114
rect 142 14 146 114
rect 264 102 268 108
rect 410 92 414 200
rect 628 138 632 295
rect 713 168 717 230
rect 781 168 785 230
rect 1057 170 1061 190
rect 1125 170 1129 295
rect 1611 277 2151 281
rect 1393 212 1397 214
rect 1395 202 1397 212
rect 903 160 907 166
rect 713 124 717 148
rect 781 124 785 148
rect 1247 162 1251 168
rect 903 134 907 140
rect 1057 126 1061 150
rect 1125 126 1129 150
rect 1247 136 1251 142
rect 903 118 907 124
rect 478 92 482 112
rect 588 96 592 102
rect 410 48 414 72
rect 478 48 482 72
rect 588 70 592 76
rect 588 54 592 60
rect 588 38 592 44
rect -270 -32 -266 -8
rect -202 -32 -198 -8
rect 214 10 218 30
rect 410 18 414 38
rect 478 16 482 38
rect -130 -18 -126 -12
rect -54 -18 -50 -6
rect -130 -34 -126 -28
rect -270 -88 -266 -42
rect -202 -88 -198 -42
rect -130 -50 -126 -44
rect -122 -90 -118 -70
rect -54 -90 -50 -28
rect 74 -30 78 -6
rect 142 -30 146 -6
rect 713 14 717 114
rect 781 14 785 114
rect 1247 120 1251 126
rect 903 102 907 108
rect 478 4 482 6
rect 214 -16 218 -10
rect 290 -16 294 -4
rect 853 10 857 30
rect 1057 16 1061 116
rect 1125 16 1129 116
rect 1247 104 1251 110
rect 1393 94 1397 202
rect 1611 140 1615 277
rect 1735 170 1739 233
rect 1803 170 1807 236
rect 2079 172 2083 192
rect 2147 172 2151 277
rect 2415 214 2419 216
rect 2417 204 2419 214
rect 1925 162 1929 168
rect 1735 126 1739 150
rect 1803 126 1807 150
rect 2269 164 2273 170
rect 1925 136 1929 142
rect 2079 128 2083 152
rect 2147 128 2151 152
rect 2269 138 2273 144
rect 1925 120 1929 126
rect 1461 94 1465 114
rect 1571 98 1575 104
rect 1393 50 1397 74
rect 1461 50 1465 74
rect 1571 72 1575 78
rect 1571 56 1575 62
rect 1571 40 1575 46
rect 214 -32 218 -26
rect 74 -86 78 -40
rect 142 -86 146 -40
rect 214 -48 218 -42
rect -270 -132 -266 -108
rect -202 -132 -198 -108
rect 222 -88 226 -68
rect 290 -88 294 -26
rect 713 -30 717 -6
rect 781 -30 785 -6
rect 1197 12 1201 32
rect 1393 20 1397 40
rect 1461 18 1465 40
rect 853 -16 857 -10
rect 929 -16 933 -4
rect 853 -32 857 -26
rect 713 -86 717 -40
rect 781 -86 785 -40
rect 853 -48 857 -42
rect -122 -114 -118 -110
rect -122 -134 -118 -124
rect -54 -134 -50 -110
rect 74 -118 78 -106
rect -16 -122 78 -118
rect 74 -130 78 -122
rect 142 -130 146 -106
rect 861 -88 865 -68
rect 929 -88 933 -26
rect 1057 -28 1061 -4
rect 1125 -28 1129 -4
rect 1735 16 1739 116
rect 1803 16 1807 116
rect 2269 122 2273 128
rect 1925 104 1929 110
rect 1461 6 1465 8
rect 1197 -14 1201 -8
rect 1273 -14 1277 -2
rect 1875 12 1879 32
rect 2079 18 2083 118
rect 2147 18 2151 118
rect 2269 106 2273 112
rect 2415 96 2419 204
rect 2633 142 2637 299
rect 2718 172 2722 235
rect 2786 172 2790 236
rect 3062 174 3066 194
rect 3130 174 3134 299
rect 3398 216 3402 218
rect 3400 206 3402 216
rect 2908 164 2912 170
rect 2718 128 2722 152
rect 2786 128 2790 152
rect 3252 166 3256 172
rect 2908 138 2912 144
rect 3062 130 3066 154
rect 3130 130 3134 154
rect 3252 140 3256 146
rect 2908 122 2912 128
rect 2483 96 2487 116
rect 2593 100 2597 106
rect 2415 52 2419 76
rect 2483 52 2487 76
rect 2593 74 2597 80
rect 2593 58 2597 64
rect 2593 42 2597 48
rect 1197 -30 1201 -24
rect 1057 -84 1061 -38
rect 1125 -84 1129 -38
rect 1197 -46 1201 -40
rect 222 -112 226 -108
rect -270 -162 -266 -142
rect -202 -162 -198 -142
rect 222 -132 226 -122
rect 290 -132 294 -108
rect 328 -120 342 -116
rect 713 -130 717 -106
rect 781 -130 785 -106
rect 1205 -86 1209 -66
rect 1273 -86 1277 -24
rect 1735 -28 1739 -4
rect 1803 -28 1807 -4
rect 2219 14 2223 34
rect 2415 22 2419 42
rect 2483 20 2487 42
rect 1875 -14 1879 -8
rect 1951 -14 1955 -2
rect 1875 -30 1879 -24
rect 1735 -84 1739 -38
rect 1803 -84 1807 -38
rect 1875 -46 1879 -40
rect 861 -112 865 -108
rect -122 -164 -118 -144
rect -54 -164 -50 -144
rect 74 -160 78 -140
rect 142 -160 146 -140
rect 861 -132 865 -122
rect 929 -132 933 -108
rect 1057 -116 1061 -104
rect 967 -120 1061 -116
rect 1057 -128 1061 -120
rect 1125 -128 1129 -104
rect 1883 -86 1887 -66
rect 1951 -86 1955 -24
rect 2079 -26 2083 -2
rect 2147 -26 2151 -2
rect 2718 18 2722 118
rect 2786 18 2790 118
rect 3252 124 3256 130
rect 2908 106 2912 112
rect 2483 8 2487 10
rect 2219 -12 2223 -6
rect 2295 -12 2299 0
rect 2858 14 2862 34
rect 3062 20 3066 120
rect 3130 20 3134 120
rect 3252 108 3256 114
rect 3398 98 3402 206
rect 3616 144 3620 181
rect 3466 98 3470 118
rect 3576 102 3580 108
rect 3398 54 3402 78
rect 3466 54 3470 78
rect 3576 76 3580 82
rect 3576 60 3580 66
rect 3576 44 3580 50
rect 2219 -28 2223 -22
rect 2079 -82 2083 -36
rect 2147 -82 2151 -36
rect 2219 -44 2223 -38
rect 1205 -110 1209 -106
rect 222 -162 226 -142
rect 290 -162 294 -142
rect 713 -160 717 -140
rect 781 -160 785 -140
rect 1205 -130 1209 -120
rect 1273 -130 1277 -106
rect 1311 -118 1325 -114
rect 1735 -128 1739 -104
rect 1803 -128 1807 -104
rect 2227 -84 2231 -64
rect 2295 -84 2299 -22
rect 2718 -26 2722 -2
rect 2786 -26 2790 -2
rect 3202 16 3206 36
rect 3398 24 3402 44
rect 3466 22 3470 44
rect 2858 -12 2862 -6
rect 2934 -12 2938 0
rect 2858 -28 2862 -22
rect 2718 -82 2722 -36
rect 2786 -82 2790 -36
rect 2858 -44 2862 -38
rect 1883 -110 1887 -106
rect 861 -162 865 -142
rect 929 -162 933 -142
rect 1057 -158 1061 -138
rect 1125 -158 1129 -138
rect 1883 -130 1887 -120
rect 1951 -130 1955 -106
rect 2079 -114 2083 -102
rect 1989 -118 2083 -114
rect 2079 -126 2083 -118
rect 2147 -126 2151 -102
rect 2866 -84 2870 -64
rect 2934 -84 2938 -22
rect 3062 -24 3066 0
rect 3130 -24 3134 0
rect 3466 10 3470 12
rect 3202 -10 3206 -4
rect 3278 -10 3282 2
rect 3202 -26 3206 -20
rect 3062 -80 3066 -34
rect 3130 -80 3134 -34
rect 3202 -42 3206 -36
rect 2227 -108 2231 -104
rect 1205 -160 1209 -140
rect 1273 -160 1277 -140
rect 1735 -158 1739 -138
rect 1803 -158 1807 -138
rect 2227 -128 2231 -118
rect 2295 -128 2299 -104
rect 2333 -116 2348 -112
rect 2718 -126 2722 -102
rect 2786 -126 2790 -102
rect 3210 -82 3214 -62
rect 3278 -82 3282 -20
rect 2866 -108 2870 -104
rect 1883 -160 1887 -140
rect 1951 -160 1955 -140
rect 2079 -156 2083 -136
rect 2147 -156 2151 -136
rect 2866 -128 2870 -118
rect 2934 -128 2938 -104
rect 3062 -112 3066 -100
rect 2972 -116 3066 -112
rect 3062 -124 3066 -116
rect 3130 -124 3134 -100
rect 3210 -106 3214 -102
rect 2227 -158 2231 -138
rect 2295 -158 2299 -138
rect 2718 -156 2722 -136
rect 2786 -156 2790 -136
rect 3210 -126 3214 -116
rect 3278 -126 3282 -102
rect 3316 -114 3331 -110
rect 2866 -158 2870 -138
rect 2934 -158 2938 -138
rect 3062 -154 3066 -134
rect 3130 -154 3134 -134
rect 3210 -156 3214 -136
rect 3278 -156 3282 -136
<< ndiffusion >>
rect -288 112 -286 122
rect -276 112 -270 122
rect -266 112 -202 122
rect -198 112 -194 122
rect -184 112 -182 122
rect -102 106 -100 116
rect -90 106 -80 116
rect -76 106 -66 116
rect -56 106 -54 116
rect 56 114 58 124
rect 68 114 74 124
rect 78 114 142 124
rect 146 114 150 124
rect 160 114 162 124
rect 242 108 244 118
rect 254 108 264 118
rect 268 108 278 118
rect 288 108 290 118
rect 695 114 697 124
rect 707 114 713 124
rect 717 114 781 124
rect 785 114 789 124
rect 799 114 801 124
rect 392 38 394 48
rect 404 38 410 48
rect 414 38 436 48
rect 446 38 478 48
rect 482 38 486 48
rect 496 38 498 48
rect 566 44 568 54
rect 578 44 588 54
rect 592 44 602 54
rect 612 44 614 54
rect -288 -42 -286 -32
rect -276 -42 -270 -32
rect -266 -42 -202 -32
rect -198 -42 -194 -32
rect -184 -42 -182 -32
rect -152 -44 -150 -34
rect -140 -44 -130 -34
rect -126 -44 -116 -34
rect -106 -44 -104 -34
rect 881 108 883 118
rect 893 108 903 118
rect 907 108 917 118
rect 927 108 929 118
rect 1039 116 1041 126
rect 1051 116 1057 126
rect 1061 116 1125 126
rect 1129 116 1133 126
rect 1143 116 1145 126
rect 1225 110 1227 120
rect 1237 110 1247 120
rect 1251 110 1261 120
rect 1271 110 1273 120
rect 1717 116 1719 126
rect 1729 116 1735 126
rect 1739 116 1803 126
rect 1807 116 1811 126
rect 1821 116 1823 126
rect 1375 40 1377 50
rect 1387 40 1393 50
rect 1397 40 1419 50
rect 1429 40 1461 50
rect 1465 40 1469 50
rect 1479 40 1481 50
rect 1549 46 1551 56
rect 1561 46 1571 56
rect 1575 46 1585 56
rect 1595 46 1597 56
rect 56 -40 58 -30
rect 68 -40 74 -30
rect 78 -40 142 -30
rect 146 -40 150 -30
rect 160 -40 162 -30
rect 192 -42 194 -32
rect 204 -42 214 -32
rect 218 -42 228 -32
rect 238 -42 240 -32
rect 695 -40 697 -30
rect 707 -40 713 -30
rect 717 -40 781 -30
rect 785 -40 789 -30
rect 799 -40 801 -30
rect 831 -42 833 -32
rect 843 -42 853 -32
rect 857 -42 867 -32
rect 877 -42 879 -32
rect -288 -142 -286 -132
rect -276 -142 -270 -132
rect -266 -142 -244 -132
rect -234 -142 -202 -132
rect -198 -142 -194 -132
rect -184 -142 -182 -132
rect 1903 110 1905 120
rect 1915 110 1925 120
rect 1929 110 1939 120
rect 1949 110 1951 120
rect 2061 118 2063 128
rect 2073 118 2079 128
rect 2083 118 2147 128
rect 2151 118 2155 128
rect 2165 118 2167 128
rect 2247 112 2249 122
rect 2259 112 2269 122
rect 2273 112 2283 122
rect 2293 112 2295 122
rect 2700 118 2702 128
rect 2712 118 2718 128
rect 2722 118 2786 128
rect 2790 118 2794 128
rect 2804 118 2806 128
rect 2397 42 2399 52
rect 2409 42 2415 52
rect 2419 42 2441 52
rect 2451 42 2483 52
rect 2487 42 2491 52
rect 2501 42 2503 52
rect 2571 48 2573 58
rect 2583 48 2593 58
rect 2597 48 2607 58
rect 2617 48 2619 58
rect 1039 -38 1041 -28
rect 1051 -38 1057 -28
rect 1061 -38 1125 -28
rect 1129 -38 1133 -28
rect 1143 -38 1145 -28
rect 1175 -40 1177 -30
rect 1187 -40 1197 -30
rect 1201 -40 1211 -30
rect 1221 -40 1223 -30
rect -140 -144 -138 -134
rect -128 -144 -122 -134
rect -118 -144 -96 -134
rect -86 -144 -54 -134
rect -50 -144 -46 -134
rect -36 -144 -34 -134
rect 56 -140 58 -130
rect 68 -140 74 -130
rect 78 -140 100 -130
rect 110 -140 142 -130
rect 146 -140 150 -130
rect 160 -140 162 -130
rect 1717 -38 1719 -28
rect 1729 -38 1735 -28
rect 1739 -38 1803 -28
rect 1807 -38 1811 -28
rect 1821 -38 1823 -28
rect 1853 -40 1855 -30
rect 1865 -40 1875 -30
rect 1879 -40 1889 -30
rect 1899 -40 1901 -30
rect 204 -142 206 -132
rect 216 -142 222 -132
rect 226 -142 248 -132
rect 258 -142 290 -132
rect 294 -142 298 -132
rect 308 -142 310 -132
rect 695 -140 697 -130
rect 707 -140 713 -130
rect 717 -140 739 -130
rect 749 -140 781 -130
rect 785 -140 789 -130
rect 799 -140 801 -130
rect 2886 112 2888 122
rect 2898 112 2908 122
rect 2912 112 2922 122
rect 2932 112 2934 122
rect 3044 120 3046 130
rect 3056 120 3062 130
rect 3066 120 3130 130
rect 3134 120 3138 130
rect 3148 120 3150 130
rect 3230 114 3232 124
rect 3242 114 3252 124
rect 3256 114 3266 124
rect 3276 114 3278 124
rect 3380 44 3382 54
rect 3392 44 3398 54
rect 3402 44 3424 54
rect 3434 44 3466 54
rect 3470 44 3474 54
rect 3484 44 3486 54
rect 3554 50 3556 60
rect 3566 50 3576 60
rect 3580 50 3590 60
rect 3600 50 3602 60
rect 2061 -36 2063 -26
rect 2073 -36 2079 -26
rect 2083 -36 2147 -26
rect 2151 -36 2155 -26
rect 2165 -36 2167 -26
rect 2197 -38 2199 -28
rect 2209 -38 2219 -28
rect 2223 -38 2233 -28
rect 2243 -38 2245 -28
rect 843 -142 845 -132
rect 855 -142 861 -132
rect 865 -142 887 -132
rect 897 -142 929 -132
rect 933 -142 937 -132
rect 947 -142 949 -132
rect 1039 -138 1041 -128
rect 1051 -138 1057 -128
rect 1061 -138 1083 -128
rect 1093 -138 1125 -128
rect 1129 -138 1133 -128
rect 1143 -138 1145 -128
rect 2700 -36 2702 -26
rect 2712 -36 2718 -26
rect 2722 -36 2786 -26
rect 2790 -36 2794 -26
rect 2804 -36 2806 -26
rect 2836 -38 2838 -28
rect 2848 -38 2858 -28
rect 2862 -38 2872 -28
rect 2882 -38 2884 -28
rect 1187 -140 1189 -130
rect 1199 -140 1205 -130
rect 1209 -140 1231 -130
rect 1241 -140 1273 -130
rect 1277 -140 1281 -130
rect 1291 -140 1293 -130
rect 1717 -138 1719 -128
rect 1729 -138 1735 -128
rect 1739 -138 1761 -128
rect 1771 -138 1803 -128
rect 1807 -138 1811 -128
rect 1821 -138 1823 -128
rect 3044 -34 3046 -24
rect 3056 -34 3062 -24
rect 3066 -34 3130 -24
rect 3134 -34 3138 -24
rect 3148 -34 3150 -24
rect 3180 -36 3182 -26
rect 3192 -36 3202 -26
rect 3206 -36 3216 -26
rect 3226 -36 3228 -26
rect 1865 -140 1867 -130
rect 1877 -140 1883 -130
rect 1887 -140 1909 -130
rect 1919 -140 1951 -130
rect 1955 -140 1959 -130
rect 1969 -140 1971 -130
rect 2061 -136 2063 -126
rect 2073 -136 2079 -126
rect 2083 -136 2105 -126
rect 2115 -136 2147 -126
rect 2151 -136 2155 -126
rect 2165 -136 2167 -126
rect 2209 -138 2211 -128
rect 2221 -138 2227 -128
rect 2231 -138 2253 -128
rect 2263 -138 2295 -128
rect 2299 -138 2303 -128
rect 2313 -138 2315 -128
rect 2700 -136 2702 -126
rect 2712 -136 2718 -126
rect 2722 -136 2744 -126
rect 2754 -136 2786 -126
rect 2790 -136 2794 -126
rect 2804 -136 2806 -126
rect 2848 -138 2850 -128
rect 2860 -138 2866 -128
rect 2870 -138 2892 -128
rect 2902 -138 2934 -128
rect 2938 -138 2942 -128
rect 2952 -138 2954 -128
rect 3044 -134 3046 -124
rect 3056 -134 3062 -124
rect 3066 -134 3088 -124
rect 3098 -134 3130 -124
rect 3134 -134 3138 -124
rect 3148 -134 3150 -124
rect 3192 -136 3194 -126
rect 3204 -136 3210 -126
rect 3214 -136 3236 -126
rect 3246 -136 3278 -126
rect 3282 -136 3286 -126
rect 3296 -136 3298 -126
<< pdiffusion >>
rect -288 160 -270 166
rect -288 150 -286 160
rect -276 150 -270 160
rect -288 146 -270 150
rect -266 160 -202 166
rect -266 150 -244 160
rect -234 150 -202 160
rect -266 146 -202 150
rect -198 160 -182 166
rect -198 150 -194 160
rect -184 150 -182 160
rect 56 162 74 168
rect -198 146 -182 150
rect -102 154 -80 158
rect -102 144 -100 154
rect -90 144 -80 154
rect -102 138 -80 144
rect -76 154 -54 158
rect -76 144 -66 154
rect -56 144 -54 154
rect 56 152 58 162
rect 68 152 74 162
rect 56 148 74 152
rect 78 162 142 168
rect 78 152 100 162
rect 110 152 142 162
rect 78 148 142 152
rect 146 162 162 168
rect 146 152 150 162
rect 160 152 162 162
rect 146 148 162 152
rect 242 156 264 160
rect -76 138 -54 144
rect 242 146 244 156
rect 254 146 264 156
rect 242 140 264 146
rect 268 156 290 160
rect 268 146 278 156
rect 288 146 290 156
rect 268 140 290 146
rect -288 6 -270 12
rect -288 -4 -286 6
rect -276 -4 -270 6
rect -288 -8 -270 -4
rect -266 6 -202 12
rect -266 -4 -244 6
rect -234 -4 -202 6
rect -266 -8 -202 -4
rect -198 6 -182 12
rect 695 162 713 168
rect 695 152 697 162
rect 707 152 713 162
rect 695 148 713 152
rect 717 162 781 168
rect 717 152 739 162
rect 749 152 781 162
rect 717 148 781 152
rect 785 162 801 168
rect 785 152 789 162
rect 799 152 801 162
rect 1039 164 1057 170
rect 785 148 801 152
rect 881 156 903 160
rect 881 146 883 156
rect 893 146 903 156
rect 881 140 903 146
rect 907 156 929 160
rect 907 146 917 156
rect 927 146 929 156
rect 1039 154 1041 164
rect 1051 154 1057 164
rect 1039 150 1057 154
rect 1061 164 1125 170
rect 1061 154 1083 164
rect 1093 154 1125 164
rect 1061 150 1125 154
rect 1129 164 1145 170
rect 1129 154 1133 164
rect 1143 154 1145 164
rect 1129 150 1145 154
rect 1225 158 1247 162
rect 907 140 929 146
rect 1225 148 1227 158
rect 1237 148 1247 158
rect 1225 142 1247 148
rect 1251 158 1273 162
rect 1251 148 1261 158
rect 1271 148 1273 158
rect 1251 142 1273 148
rect 566 92 588 96
rect 392 86 410 92
rect 392 76 394 86
rect 404 76 410 86
rect 392 72 410 76
rect 414 72 478 92
rect 482 86 498 92
rect 482 76 486 86
rect 496 76 498 86
rect 566 82 568 92
rect 578 82 588 92
rect 566 76 588 82
rect 592 92 614 96
rect 592 82 602 92
rect 612 82 614 92
rect 592 76 614 82
rect 482 72 498 76
rect 56 8 74 14
rect -198 -4 -194 6
rect -184 -4 -182 6
rect -198 -8 -182 -4
rect -152 4 -130 8
rect -152 -6 -150 4
rect -140 -6 -130 4
rect -152 -12 -130 -6
rect -126 4 -104 8
rect -126 -6 -116 4
rect -106 -6 -104 4
rect 56 -2 58 8
rect 68 -2 74 8
rect 56 -6 74 -2
rect 78 8 142 14
rect 78 -2 100 8
rect 110 -2 142 8
rect 78 -6 142 -2
rect 146 8 162 14
rect 146 -2 150 8
rect 160 -2 162 8
rect 146 -6 162 -2
rect 192 6 214 10
rect 192 -4 194 6
rect 204 -4 214 6
rect -126 -12 -104 -6
rect -288 -94 -270 -88
rect -288 -104 -286 -94
rect -276 -104 -270 -94
rect -288 -108 -270 -104
rect -266 -108 -202 -88
rect -198 -94 -182 -88
rect 192 -10 214 -4
rect 218 6 240 10
rect 218 -4 228 6
rect 238 -4 240 6
rect 695 8 713 14
rect 695 -2 697 8
rect 707 -2 713 8
rect 218 -10 240 -4
rect 695 -6 713 -2
rect 717 8 781 14
rect 717 -2 739 8
rect 749 -2 781 8
rect 717 -6 781 -2
rect 785 8 801 14
rect 1717 164 1735 170
rect 1717 154 1719 164
rect 1729 154 1735 164
rect 1717 150 1735 154
rect 1739 164 1803 170
rect 1739 154 1761 164
rect 1771 154 1803 164
rect 1739 150 1803 154
rect 1807 164 1823 170
rect 1807 154 1811 164
rect 1821 154 1823 164
rect 2061 166 2079 172
rect 1807 150 1823 154
rect 1903 158 1925 162
rect 1903 148 1905 158
rect 1915 148 1925 158
rect 1903 142 1925 148
rect 1929 158 1951 162
rect 1929 148 1939 158
rect 1949 148 1951 158
rect 2061 156 2063 166
rect 2073 156 2079 166
rect 2061 152 2079 156
rect 2083 166 2147 172
rect 2083 156 2105 166
rect 2115 156 2147 166
rect 2083 152 2147 156
rect 2151 166 2167 172
rect 2151 156 2155 166
rect 2165 156 2167 166
rect 2151 152 2167 156
rect 2247 160 2269 164
rect 1929 142 1951 148
rect 2247 150 2249 160
rect 2259 150 2269 160
rect 2247 144 2269 150
rect 2273 160 2295 164
rect 2273 150 2283 160
rect 2293 150 2295 160
rect 2273 144 2295 150
rect 1549 94 1571 98
rect 1375 88 1393 94
rect 1375 78 1377 88
rect 1387 78 1393 88
rect 1375 74 1393 78
rect 1397 74 1461 94
rect 1465 88 1481 94
rect 1465 78 1469 88
rect 1479 78 1481 88
rect 1549 84 1551 94
rect 1561 84 1571 94
rect 1549 78 1571 84
rect 1575 94 1597 98
rect 1575 84 1585 94
rect 1595 84 1597 94
rect 1575 78 1597 84
rect 1465 74 1481 78
rect 1039 10 1057 16
rect 785 -2 789 8
rect 799 -2 801 8
rect 785 -6 801 -2
rect 831 6 853 10
rect 831 -4 833 6
rect 843 -4 853 6
rect -198 -104 -194 -94
rect -184 -104 -182 -94
rect -198 -108 -182 -104
rect -140 -96 -122 -90
rect -140 -106 -138 -96
rect -128 -106 -122 -96
rect -140 -110 -122 -106
rect -118 -110 -54 -90
rect -50 -96 -34 -90
rect -50 -106 -46 -96
rect -36 -106 -34 -96
rect 56 -92 74 -86
rect 56 -102 58 -92
rect 68 -102 74 -92
rect 56 -106 74 -102
rect 78 -106 142 -86
rect 146 -92 162 -86
rect 831 -10 853 -4
rect 857 6 879 10
rect 857 -4 867 6
rect 877 -4 879 6
rect 1039 0 1041 10
rect 1051 0 1057 10
rect 1039 -4 1057 0
rect 1061 10 1125 16
rect 1061 0 1083 10
rect 1093 0 1125 10
rect 1061 -4 1125 0
rect 1129 10 1145 16
rect 1129 0 1133 10
rect 1143 0 1145 10
rect 1129 -4 1145 0
rect 1175 8 1197 12
rect 1175 -2 1177 8
rect 1187 -2 1197 8
rect 857 -10 879 -4
rect 146 -102 150 -92
rect 160 -102 162 -92
rect 146 -106 162 -102
rect 204 -94 222 -88
rect 204 -104 206 -94
rect 216 -104 222 -94
rect -50 -110 -34 -106
rect 204 -108 222 -104
rect 226 -108 290 -88
rect 294 -94 310 -88
rect 294 -104 298 -94
rect 308 -104 310 -94
rect 294 -108 310 -104
rect 695 -92 713 -86
rect 695 -102 697 -92
rect 707 -102 713 -92
rect 695 -106 713 -102
rect 717 -106 781 -86
rect 785 -92 801 -86
rect 1175 -8 1197 -2
rect 1201 8 1223 12
rect 1201 -2 1211 8
rect 1221 -2 1223 8
rect 1717 10 1735 16
rect 1717 0 1719 10
rect 1729 0 1735 10
rect 1201 -8 1223 -2
rect 1717 -4 1735 0
rect 1739 10 1803 16
rect 1739 0 1761 10
rect 1771 0 1803 10
rect 1739 -4 1803 0
rect 1807 10 1823 16
rect 2700 166 2718 172
rect 2700 156 2702 166
rect 2712 156 2718 166
rect 2700 152 2718 156
rect 2722 166 2786 172
rect 2722 156 2744 166
rect 2754 156 2786 166
rect 2722 152 2786 156
rect 2790 166 2806 172
rect 2790 156 2794 166
rect 2804 156 2806 166
rect 3044 168 3062 174
rect 2790 152 2806 156
rect 2886 160 2908 164
rect 2886 150 2888 160
rect 2898 150 2908 160
rect 2886 144 2908 150
rect 2912 160 2934 164
rect 2912 150 2922 160
rect 2932 150 2934 160
rect 3044 158 3046 168
rect 3056 158 3062 168
rect 3044 154 3062 158
rect 3066 168 3130 174
rect 3066 158 3088 168
rect 3098 158 3130 168
rect 3066 154 3130 158
rect 3134 168 3150 174
rect 3134 158 3138 168
rect 3148 158 3150 168
rect 3134 154 3150 158
rect 3230 162 3252 166
rect 2912 144 2934 150
rect 3230 152 3232 162
rect 3242 152 3252 162
rect 3230 146 3252 152
rect 3256 162 3278 166
rect 3256 152 3266 162
rect 3276 152 3278 162
rect 3256 146 3278 152
rect 2571 96 2593 100
rect 2397 90 2415 96
rect 2397 80 2399 90
rect 2409 80 2415 90
rect 2397 76 2415 80
rect 2419 76 2483 96
rect 2487 90 2503 96
rect 2487 80 2491 90
rect 2501 80 2503 90
rect 2571 86 2573 96
rect 2583 86 2593 96
rect 2571 80 2593 86
rect 2597 96 2619 100
rect 2597 86 2607 96
rect 2617 86 2619 96
rect 2597 80 2619 86
rect 2487 76 2503 80
rect 2061 12 2079 18
rect 1807 0 1811 10
rect 1821 0 1823 10
rect 1807 -4 1823 0
rect 1853 8 1875 12
rect 1853 -2 1855 8
rect 1865 -2 1875 8
rect 785 -102 789 -92
rect 799 -102 801 -92
rect 785 -106 801 -102
rect 843 -94 861 -88
rect 843 -104 845 -94
rect 855 -104 861 -94
rect 843 -108 861 -104
rect 865 -108 929 -88
rect 933 -94 949 -88
rect 933 -104 937 -94
rect 947 -104 949 -94
rect 1039 -90 1057 -84
rect 1039 -100 1041 -90
rect 1051 -100 1057 -90
rect 1039 -104 1057 -100
rect 1061 -104 1125 -84
rect 1129 -90 1145 -84
rect 1853 -8 1875 -2
rect 1879 8 1901 12
rect 1879 -2 1889 8
rect 1899 -2 1901 8
rect 2061 2 2063 12
rect 2073 2 2079 12
rect 2061 -2 2079 2
rect 2083 12 2147 18
rect 2083 2 2105 12
rect 2115 2 2147 12
rect 2083 -2 2147 2
rect 2151 12 2167 18
rect 2151 2 2155 12
rect 2165 2 2167 12
rect 2151 -2 2167 2
rect 2197 10 2219 14
rect 2197 0 2199 10
rect 2209 0 2219 10
rect 1879 -8 1901 -2
rect 1129 -100 1133 -90
rect 1143 -100 1145 -90
rect 1129 -104 1145 -100
rect 1187 -92 1205 -86
rect 1187 -102 1189 -92
rect 1199 -102 1205 -92
rect 933 -108 949 -104
rect 1187 -106 1205 -102
rect 1209 -106 1273 -86
rect 1277 -92 1293 -86
rect 1277 -102 1281 -92
rect 1291 -102 1293 -92
rect 1277 -106 1293 -102
rect 1717 -90 1735 -84
rect 1717 -100 1719 -90
rect 1729 -100 1735 -90
rect 1717 -104 1735 -100
rect 1739 -104 1803 -84
rect 1807 -90 1823 -84
rect 2197 -6 2219 0
rect 2223 10 2245 14
rect 2223 0 2233 10
rect 2243 0 2245 10
rect 2700 12 2718 18
rect 2700 2 2702 12
rect 2712 2 2718 12
rect 2223 -6 2245 0
rect 2700 -2 2718 2
rect 2722 12 2786 18
rect 2722 2 2744 12
rect 2754 2 2786 12
rect 2722 -2 2786 2
rect 2790 12 2806 18
rect 3554 98 3576 102
rect 3380 92 3398 98
rect 3380 82 3382 92
rect 3392 82 3398 92
rect 3380 78 3398 82
rect 3402 78 3466 98
rect 3470 92 3486 98
rect 3470 82 3474 92
rect 3484 82 3486 92
rect 3554 88 3556 98
rect 3566 88 3576 98
rect 3554 82 3576 88
rect 3580 98 3602 102
rect 3580 88 3590 98
rect 3600 88 3602 98
rect 3580 82 3602 88
rect 3470 78 3486 82
rect 3044 14 3062 20
rect 2790 2 2794 12
rect 2804 2 2806 12
rect 2790 -2 2806 2
rect 2836 10 2858 14
rect 2836 0 2838 10
rect 2848 0 2858 10
rect 1807 -100 1811 -90
rect 1821 -100 1823 -90
rect 1807 -104 1823 -100
rect 1865 -92 1883 -86
rect 1865 -102 1867 -92
rect 1877 -102 1883 -92
rect 1865 -106 1883 -102
rect 1887 -106 1951 -86
rect 1955 -92 1971 -86
rect 1955 -102 1959 -92
rect 1969 -102 1971 -92
rect 2061 -88 2079 -82
rect 2061 -98 2063 -88
rect 2073 -98 2079 -88
rect 2061 -102 2079 -98
rect 2083 -102 2147 -82
rect 2151 -88 2167 -82
rect 2836 -6 2858 0
rect 2862 10 2884 14
rect 2862 0 2872 10
rect 2882 0 2884 10
rect 3044 4 3046 14
rect 3056 4 3062 14
rect 3044 0 3062 4
rect 3066 14 3130 20
rect 3066 4 3088 14
rect 3098 4 3130 14
rect 3066 0 3130 4
rect 3134 14 3150 20
rect 3134 4 3138 14
rect 3148 4 3150 14
rect 3134 0 3150 4
rect 3180 12 3202 16
rect 3180 2 3182 12
rect 3192 2 3202 12
rect 2862 -6 2884 0
rect 2151 -98 2155 -88
rect 2165 -98 2167 -88
rect 2151 -102 2167 -98
rect 2209 -90 2227 -84
rect 2209 -100 2211 -90
rect 2221 -100 2227 -90
rect 1955 -106 1971 -102
rect 2209 -104 2227 -100
rect 2231 -104 2295 -84
rect 2299 -90 2315 -84
rect 2299 -100 2303 -90
rect 2313 -100 2315 -90
rect 2299 -104 2315 -100
rect 2700 -88 2718 -82
rect 2700 -98 2702 -88
rect 2712 -98 2718 -88
rect 2700 -102 2718 -98
rect 2722 -102 2786 -82
rect 2790 -88 2806 -82
rect 3180 -4 3202 2
rect 3206 12 3228 16
rect 3206 2 3216 12
rect 3226 2 3228 12
rect 3206 -4 3228 2
rect 2790 -98 2794 -88
rect 2804 -98 2806 -88
rect 2790 -102 2806 -98
rect 2848 -90 2866 -84
rect 2848 -100 2850 -90
rect 2860 -100 2866 -90
rect 2848 -104 2866 -100
rect 2870 -104 2934 -84
rect 2938 -90 2954 -84
rect 2938 -100 2942 -90
rect 2952 -100 2954 -90
rect 3044 -86 3062 -80
rect 3044 -96 3046 -86
rect 3056 -96 3062 -86
rect 3044 -100 3062 -96
rect 3066 -100 3130 -80
rect 3134 -86 3150 -80
rect 3134 -96 3138 -86
rect 3148 -96 3150 -86
rect 3134 -100 3150 -96
rect 3192 -88 3210 -82
rect 3192 -98 3194 -88
rect 3204 -98 3210 -88
rect 2938 -104 2954 -100
rect 3192 -102 3210 -98
rect 3214 -102 3278 -82
rect 3282 -88 3298 -82
rect 3282 -98 3286 -88
rect 3296 -98 3298 -88
rect 3282 -102 3298 -98
<< metal1 >>
rect 336 200 402 210
rect 1319 202 1385 212
rect 2341 204 2407 214
rect 3324 206 3390 216
rect 2964 184 3318 186
rect 1981 182 3318 184
rect 959 180 3318 182
rect -24 178 3318 180
rect -298 176 3318 178
rect -298 174 2974 176
rect -298 172 1991 174
rect -298 170 969 172
rect -298 168 -14 170
rect -286 160 -276 168
rect -194 160 -184 168
rect -100 154 -90 168
rect -244 140 -234 150
rect -244 132 -164 140
rect -66 132 -56 144
rect -244 130 -86 132
rect -194 122 -184 130
rect -174 122 -86 130
rect -66 122 -48 132
rect -66 116 -56 122
rect -286 106 -276 112
rect -310 100 -164 106
rect -100 100 -90 106
rect -310 96 -90 100
rect -310 -48 -300 96
rect -174 90 -90 96
rect -24 24 -14 168
rect 58 162 68 170
rect 150 162 160 170
rect 244 156 254 170
rect 100 142 110 152
rect 100 134 180 142
rect 278 134 288 146
rect 100 132 258 134
rect 150 124 160 132
rect 170 124 258 132
rect 278 124 296 134
rect 278 118 288 124
rect 58 108 68 114
rect -286 14 -14 24
rect -286 6 -276 14
rect -194 6 -184 14
rect -150 12 -14 14
rect -150 4 -140 12
rect -244 -14 -234 -4
rect -244 -18 -164 -14
rect -116 -18 -106 -6
rect -244 -24 -136 -18
rect -194 -32 -184 -24
rect -174 -28 -136 -24
rect -116 -28 -60 -18
rect -116 -34 -106 -28
rect -286 -48 -276 -42
rect -150 -48 -140 -44
rect -310 -58 -140 -48
rect -310 -150 -300 -58
rect -24 -76 -14 12
rect -286 -86 -14 -76
rect 34 102 180 108
rect 244 102 254 108
rect 34 98 254 102
rect 34 -46 44 98
rect 170 92 254 98
rect 320 104 330 170
rect 697 162 707 170
rect 789 162 799 170
rect 883 156 893 170
rect 739 142 749 152
rect 739 134 819 142
rect 917 134 927 146
rect 739 132 897 134
rect 394 104 578 106
rect 392 96 578 104
rect 392 94 404 96
rect 320 26 330 94
rect 394 86 404 94
rect 568 92 578 96
rect 486 66 496 76
rect 602 70 612 82
rect 624 70 634 128
rect 789 124 799 132
rect 809 124 897 132
rect 917 124 935 134
rect 917 118 927 124
rect 697 108 707 114
rect 506 66 582 70
rect 436 60 582 66
rect 602 60 634 70
rect 673 102 819 108
rect 883 102 893 108
rect 673 98 893 102
rect 436 56 516 60
rect 436 48 446 56
rect 602 54 612 60
rect 58 16 330 26
rect 58 8 68 16
rect 150 8 160 16
rect 194 14 330 16
rect 194 6 204 14
rect 100 -12 110 -2
rect 100 -16 180 -12
rect 228 -16 238 -4
rect 100 -22 208 -16
rect 150 -30 160 -22
rect 170 -26 208 -22
rect 228 -26 284 -16
rect 228 -32 238 -26
rect 58 -46 68 -40
rect 194 -46 204 -42
rect 34 -56 204 -46
rect -286 -94 -276 -86
rect -194 -114 -184 -104
rect -138 -96 -128 -86
rect -244 -124 -128 -114
rect -46 -116 -36 -106
rect -244 -132 -234 -124
rect -96 -126 -26 -116
rect -96 -134 -86 -126
rect -286 -150 -276 -142
rect -194 -150 -184 -142
rect -138 -150 -128 -144
rect -46 -150 -36 -144
rect 34 -148 44 -56
rect 320 -74 330 14
rect 58 -84 330 -74
rect 394 32 404 38
rect 486 32 496 38
rect 568 32 578 44
rect 394 22 578 32
rect 58 -92 68 -84
rect 150 -112 160 -102
rect 206 -94 216 -84
rect 100 -122 216 -112
rect 298 -114 308 -104
rect 100 -130 110 -122
rect 248 -124 318 -114
rect 248 -132 258 -124
rect 58 -148 68 -140
rect 150 -148 160 -140
rect 206 -148 216 -142
rect 298 -148 308 -142
rect 394 -148 404 22
rect 516 20 578 22
rect 454 6 472 16
rect 673 -46 683 98
rect 809 92 893 98
rect 959 26 969 170
rect 1041 164 1051 172
rect 1133 164 1143 172
rect 1227 158 1237 172
rect 1083 144 1093 154
rect 1083 136 1163 144
rect 1261 136 1271 148
rect 1083 134 1241 136
rect 1133 126 1143 134
rect 1153 126 1241 134
rect 1261 126 1279 136
rect 1261 120 1271 126
rect 1041 110 1051 116
rect 697 16 969 26
rect 697 8 707 16
rect 789 8 799 16
rect 833 14 969 16
rect 833 6 843 14
rect 739 -12 749 -2
rect 739 -16 819 -12
rect 867 -16 877 -4
rect 739 -22 847 -16
rect 789 -30 799 -22
rect 809 -26 847 -22
rect 867 -26 923 -16
rect 867 -32 877 -26
rect 697 -46 707 -40
rect 833 -46 843 -42
rect 673 -56 843 -46
rect 673 -148 683 -56
rect 959 -74 969 14
rect 697 -84 969 -74
rect 1017 104 1163 110
rect 1227 104 1237 110
rect 1017 100 1237 104
rect 1017 -44 1027 100
rect 1153 94 1237 100
rect 1303 106 1313 172
rect 1719 164 1729 172
rect 1811 164 1821 172
rect 1905 158 1915 172
rect 1761 144 1771 154
rect 1761 136 1841 144
rect 1939 136 1949 148
rect 1761 134 1919 136
rect 1377 106 1561 108
rect 1375 98 1561 106
rect 1375 96 1387 98
rect 1303 28 1313 96
rect 1377 88 1387 96
rect 1551 94 1561 98
rect 1469 68 1479 78
rect 1585 72 1595 84
rect 1607 72 1617 130
rect 1811 126 1821 134
rect 1831 126 1919 134
rect 1939 126 1957 136
rect 1939 120 1949 126
rect 1719 110 1729 116
rect 1489 68 1565 72
rect 1419 62 1565 68
rect 1585 62 1617 72
rect 1695 104 1841 110
rect 1905 104 1915 110
rect 1695 100 1915 104
rect 1419 58 1499 62
rect 1419 50 1429 58
rect 1585 56 1595 62
rect 1041 18 1313 28
rect 1041 10 1051 18
rect 1133 10 1143 18
rect 1177 16 1313 18
rect 1177 8 1187 16
rect 1083 -10 1093 0
rect 1083 -14 1163 -10
rect 1211 -14 1221 -2
rect 1083 -20 1191 -14
rect 1133 -28 1143 -20
rect 1153 -24 1191 -20
rect 1211 -24 1267 -14
rect 1211 -30 1221 -24
rect 1041 -44 1051 -38
rect 1177 -44 1187 -40
rect 1017 -54 1187 -44
rect 697 -92 707 -84
rect 789 -112 799 -102
rect 845 -94 855 -84
rect 739 -122 855 -112
rect 937 -114 947 -104
rect 739 -130 749 -122
rect 887 -124 957 -114
rect 887 -132 897 -124
rect 697 -148 707 -140
rect 789 -148 799 -140
rect 845 -148 855 -142
rect 937 -148 947 -142
rect 1017 -146 1027 -54
rect 1303 -72 1313 16
rect 1041 -82 1313 -72
rect 1377 34 1387 40
rect 1469 34 1479 40
rect 1551 34 1561 46
rect 1377 24 1561 34
rect 1041 -90 1051 -82
rect 1133 -110 1143 -100
rect 1189 -92 1199 -82
rect 1083 -120 1199 -110
rect 1281 -112 1291 -102
rect 1083 -128 1093 -120
rect 1231 -122 1301 -112
rect 1231 -130 1241 -122
rect 1041 -146 1051 -138
rect 1133 -146 1143 -138
rect 1189 -146 1199 -140
rect 1281 -146 1291 -140
rect 1377 -146 1387 24
rect 1499 22 1561 24
rect 1437 8 1455 18
rect 1695 -44 1705 100
rect 1831 94 1915 100
rect 1981 28 1991 172
rect 2063 166 2073 174
rect 2155 166 2165 174
rect 2249 160 2259 174
rect 2105 146 2115 156
rect 2105 138 2185 146
rect 2283 138 2293 150
rect 2105 136 2263 138
rect 2155 128 2165 136
rect 2175 128 2263 136
rect 2283 128 2301 138
rect 2283 122 2293 128
rect 2063 112 2073 118
rect 1719 18 1991 28
rect 1719 10 1729 18
rect 1811 10 1821 18
rect 1855 16 1991 18
rect 1855 8 1865 16
rect 1761 -10 1771 0
rect 1761 -14 1841 -10
rect 1889 -14 1899 -2
rect 1761 -20 1869 -14
rect 1811 -28 1821 -20
rect 1831 -24 1869 -20
rect 1889 -24 1945 -14
rect 1889 -30 1899 -24
rect 1719 -44 1729 -38
rect 1855 -44 1865 -40
rect 1695 -54 1865 -44
rect 1695 -145 1705 -54
rect 1981 -72 1991 16
rect 1719 -82 1991 -72
rect 2039 106 2185 112
rect 2249 106 2259 112
rect 2039 102 2259 106
rect 2039 -42 2049 102
rect 2175 96 2259 102
rect 2325 108 2335 174
rect 2702 166 2712 174
rect 2794 166 2804 174
rect 2888 160 2898 174
rect 2744 146 2754 156
rect 2744 138 2824 146
rect 2922 138 2932 150
rect 2744 136 2902 138
rect 2399 108 2583 110
rect 2397 100 2583 108
rect 2397 98 2409 100
rect 2325 30 2335 98
rect 2399 90 2409 98
rect 2573 96 2583 100
rect 2491 70 2501 80
rect 2607 74 2617 86
rect 2629 74 2639 132
rect 2794 128 2804 136
rect 2814 128 2902 136
rect 2922 128 2940 138
rect 2922 122 2932 128
rect 2702 112 2712 118
rect 2511 70 2587 74
rect 2441 64 2587 70
rect 2607 64 2639 74
rect 2678 106 2824 112
rect 2888 106 2898 112
rect 2678 102 2898 106
rect 2441 60 2521 64
rect 2441 52 2451 60
rect 2607 58 2617 64
rect 2063 20 2335 30
rect 2063 12 2073 20
rect 2155 12 2165 20
rect 2199 18 2335 20
rect 2199 10 2209 18
rect 2105 -8 2115 2
rect 2105 -12 2185 -8
rect 2233 -12 2243 0
rect 2105 -18 2213 -12
rect 2155 -26 2165 -18
rect 2175 -22 2213 -18
rect 2233 -22 2289 -12
rect 2233 -28 2243 -22
rect 2063 -42 2073 -36
rect 2199 -42 2209 -38
rect 2039 -52 2209 -42
rect 1719 -90 1729 -82
rect 1811 -110 1821 -100
rect 1867 -92 1877 -82
rect 1761 -120 1877 -110
rect 1959 -112 1969 -102
rect 1761 -128 1771 -120
rect 1909 -122 1979 -112
rect 1694 -146 1705 -145
rect 1909 -130 1919 -122
rect 1719 -146 1729 -138
rect 1811 -146 1821 -138
rect 1867 -146 1877 -140
rect 1959 -146 1969 -140
rect 2039 -144 2049 -52
rect 2325 -70 2335 18
rect 2063 -80 2335 -70
rect 2399 36 2409 42
rect 2491 36 2501 42
rect 2573 36 2583 48
rect 2399 26 2583 36
rect 2063 -88 2073 -80
rect 2155 -108 2165 -98
rect 2211 -90 2221 -80
rect 2105 -118 2221 -108
rect 2303 -110 2313 -100
rect 2105 -126 2115 -118
rect 2253 -120 2323 -110
rect 2253 -128 2263 -120
rect 2063 -144 2073 -136
rect 2155 -144 2165 -136
rect 2211 -144 2221 -138
rect 2303 -144 2313 -138
rect 2399 -144 2409 26
rect 2521 24 2583 26
rect 2459 10 2477 20
rect 2678 -42 2688 102
rect 2814 96 2898 102
rect 2964 30 2974 174
rect 3046 168 3056 176
rect 3138 168 3148 176
rect 3232 162 3242 176
rect 3088 148 3098 158
rect 3088 140 3168 148
rect 3266 140 3276 152
rect 3088 138 3246 140
rect 3138 130 3148 138
rect 3158 130 3246 138
rect 3266 130 3284 140
rect 3266 124 3276 130
rect 3046 114 3056 120
rect 2702 20 2974 30
rect 2702 12 2712 20
rect 2794 12 2804 20
rect 2838 18 2974 20
rect 2838 10 2848 18
rect 2744 -8 2754 2
rect 2744 -12 2824 -8
rect 2872 -12 2882 0
rect 2744 -18 2852 -12
rect 2794 -26 2804 -18
rect 2814 -22 2852 -18
rect 2872 -22 2928 -12
rect 2872 -28 2882 -22
rect 2702 -42 2712 -36
rect 2838 -42 2848 -38
rect 2678 -52 2848 -42
rect 2678 -144 2688 -52
rect 2964 -70 2974 18
rect 2702 -80 2974 -70
rect 3022 108 3168 114
rect 3232 108 3242 114
rect 3022 104 3242 108
rect 3022 -40 3032 104
rect 3158 98 3242 104
rect 3308 110 3318 176
rect 3382 110 3566 112
rect 3380 102 3566 110
rect 3380 100 3392 102
rect 3308 32 3318 100
rect 3382 92 3392 100
rect 3556 98 3566 102
rect 3474 72 3484 82
rect 3590 76 3600 88
rect 3612 76 3622 134
rect 3494 72 3570 76
rect 3424 66 3570 72
rect 3590 66 3622 76
rect 3424 62 3504 66
rect 3424 54 3434 62
rect 3590 60 3600 66
rect 3046 22 3318 32
rect 3046 14 3056 22
rect 3138 14 3148 22
rect 3182 20 3318 22
rect 3182 12 3192 20
rect 3088 -6 3098 4
rect 3088 -10 3168 -6
rect 3216 -10 3226 2
rect 3088 -16 3196 -10
rect 3138 -24 3148 -16
rect 3158 -20 3196 -16
rect 3216 -20 3272 -10
rect 3216 -26 3226 -20
rect 3046 -40 3056 -34
rect 3182 -40 3192 -36
rect 3022 -50 3192 -40
rect 2702 -88 2712 -80
rect 2794 -108 2804 -98
rect 2850 -90 2860 -80
rect 2744 -118 2860 -108
rect 2942 -110 2952 -100
rect 2744 -126 2754 -118
rect 2892 -120 2962 -110
rect 2892 -128 2902 -120
rect 2702 -144 2712 -136
rect 2794 -144 2804 -136
rect 2850 -144 2860 -138
rect 2942 -144 2952 -138
rect 3022 -142 3032 -50
rect 3308 -68 3318 20
rect 3046 -78 3318 -68
rect 3382 38 3392 44
rect 3474 38 3484 44
rect 3556 38 3566 50
rect 3382 28 3566 38
rect 3046 -86 3056 -78
rect 3138 -106 3148 -96
rect 3194 -88 3204 -78
rect 3088 -116 3204 -106
rect 3286 -108 3296 -98
rect 3088 -124 3098 -116
rect 3236 -118 3306 -108
rect 3236 -126 3246 -118
rect 3046 -142 3056 -134
rect 3138 -142 3148 -134
rect 3194 -142 3204 -136
rect 3286 -142 3296 -136
rect 3382 -142 3392 28
rect 3504 26 3566 28
rect 3442 12 3460 22
rect 3022 -144 3392 -142
rect 2039 -146 3392 -144
rect 1017 -148 3392 -146
rect 34 -150 3392 -148
rect -310 -152 3392 -150
rect -310 -154 3032 -152
rect -310 -156 2049 -154
rect -310 -158 1027 -156
rect -310 -160 44 -158
<< metal2 >>
rect -32 200 326 210
rect 951 202 1309 212
rect 1973 204 2331 214
rect 2956 206 3314 216
rect -32 132 -22 200
rect 951 134 961 202
rect 1973 136 1983 204
rect 2956 138 2966 206
rect -38 122 -22 132
rect 945 124 961 134
rect 1967 126 1983 136
rect 2950 128 2966 138
rect 296 16 306 124
rect 330 94 382 104
rect 1279 18 1289 126
rect 1313 96 1365 106
rect 2301 20 2311 128
rect 2335 98 2387 108
rect 3284 22 3294 130
rect 3318 100 3370 110
rect 296 6 444 16
rect 472 6 482 16
rect 1279 8 1427 18
rect 1455 8 1465 18
rect 2301 10 2449 20
rect 2477 10 2487 20
rect 3284 12 3432 22
rect 3460 12 3470 22
<< ntransistor >>
rect -270 112 -266 122
rect -202 112 -198 122
rect -80 106 -76 116
rect 74 114 78 124
rect 142 114 146 124
rect 264 108 268 118
rect 713 114 717 124
rect 781 114 785 124
rect 410 38 414 48
rect 478 38 482 48
rect 588 44 592 54
rect -270 -42 -266 -32
rect -202 -42 -198 -32
rect -130 -44 -126 -34
rect 903 108 907 118
rect 1057 116 1061 126
rect 1125 116 1129 126
rect 1247 110 1251 120
rect 1735 116 1739 126
rect 1803 116 1807 126
rect 1393 40 1397 50
rect 1461 40 1465 50
rect 1571 46 1575 56
rect 74 -40 78 -30
rect 142 -40 146 -30
rect 214 -42 218 -32
rect 713 -40 717 -30
rect 781 -40 785 -30
rect 853 -42 857 -32
rect -270 -142 -266 -132
rect -202 -142 -198 -132
rect 1925 110 1929 120
rect 2079 118 2083 128
rect 2147 118 2151 128
rect 2269 112 2273 122
rect 2718 118 2722 128
rect 2786 118 2790 128
rect 2415 42 2419 52
rect 2483 42 2487 52
rect 2593 48 2597 58
rect 1057 -38 1061 -28
rect 1125 -38 1129 -28
rect 1197 -40 1201 -30
rect -122 -144 -118 -134
rect -54 -144 -50 -134
rect 74 -140 78 -130
rect 142 -140 146 -130
rect 1735 -38 1739 -28
rect 1803 -38 1807 -28
rect 1875 -40 1879 -30
rect 222 -142 226 -132
rect 290 -142 294 -132
rect 713 -140 717 -130
rect 781 -140 785 -130
rect 2908 112 2912 122
rect 3062 120 3066 130
rect 3130 120 3134 130
rect 3252 114 3256 124
rect 3398 44 3402 54
rect 3466 44 3470 54
rect 3576 50 3580 60
rect 2079 -36 2083 -26
rect 2147 -36 2151 -26
rect 2219 -38 2223 -28
rect 861 -142 865 -132
rect 929 -142 933 -132
rect 1057 -138 1061 -128
rect 1125 -138 1129 -128
rect 2718 -36 2722 -26
rect 2786 -36 2790 -26
rect 2858 -38 2862 -28
rect 1205 -140 1209 -130
rect 1273 -140 1277 -130
rect 1735 -138 1739 -128
rect 1803 -138 1807 -128
rect 3062 -34 3066 -24
rect 3130 -34 3134 -24
rect 3202 -36 3206 -26
rect 1883 -140 1887 -130
rect 1951 -140 1955 -130
rect 2079 -136 2083 -126
rect 2147 -136 2151 -126
rect 2227 -138 2231 -128
rect 2295 -138 2299 -128
rect 2718 -136 2722 -126
rect 2786 -136 2790 -126
rect 2866 -138 2870 -128
rect 2934 -138 2938 -128
rect 3062 -134 3066 -124
rect 3130 -134 3134 -124
rect 3210 -136 3214 -126
rect 3278 -136 3282 -126
<< ptransistor >>
rect -270 146 -266 166
rect -202 146 -198 166
rect -80 138 -76 158
rect 74 148 78 168
rect 142 148 146 168
rect 264 140 268 160
rect -270 -8 -266 12
rect -202 -8 -198 12
rect 713 148 717 168
rect 781 148 785 168
rect 903 140 907 160
rect 1057 150 1061 170
rect 1125 150 1129 170
rect 1247 142 1251 162
rect 410 72 414 92
rect 478 72 482 92
rect 588 76 592 96
rect -130 -12 -126 8
rect 74 -6 78 14
rect 142 -6 146 14
rect -270 -108 -266 -88
rect -202 -108 -198 -88
rect 214 -10 218 10
rect 713 -6 717 14
rect 781 -6 785 14
rect 1735 150 1739 170
rect 1803 150 1807 170
rect 1925 142 1929 162
rect 2079 152 2083 172
rect 2147 152 2151 172
rect 2269 144 2273 164
rect 1393 74 1397 94
rect 1461 74 1465 94
rect 1571 78 1575 98
rect -122 -110 -118 -90
rect -54 -110 -50 -90
rect 74 -106 78 -86
rect 142 -106 146 -86
rect 853 -10 857 10
rect 1057 -4 1061 16
rect 1125 -4 1129 16
rect 222 -108 226 -88
rect 290 -108 294 -88
rect 713 -106 717 -86
rect 781 -106 785 -86
rect 1197 -8 1201 12
rect 1735 -4 1739 16
rect 1803 -4 1807 16
rect 2718 152 2722 172
rect 2786 152 2790 172
rect 2908 144 2912 164
rect 3062 154 3066 174
rect 3130 154 3134 174
rect 3252 146 3256 166
rect 2415 76 2419 96
rect 2483 76 2487 96
rect 2593 80 2597 100
rect 861 -108 865 -88
rect 929 -108 933 -88
rect 1057 -104 1061 -84
rect 1125 -104 1129 -84
rect 1875 -8 1879 12
rect 2079 -2 2083 18
rect 2147 -2 2151 18
rect 1205 -106 1209 -86
rect 1273 -106 1277 -86
rect 1735 -104 1739 -84
rect 1803 -104 1807 -84
rect 2219 -6 2223 14
rect 2718 -2 2722 18
rect 2786 -2 2790 18
rect 3398 78 3402 98
rect 3466 78 3470 98
rect 3576 82 3580 102
rect 1883 -106 1887 -86
rect 1951 -106 1955 -86
rect 2079 -102 2083 -82
rect 2147 -102 2151 -82
rect 2858 -6 2862 14
rect 3062 0 3066 20
rect 3130 0 3134 20
rect 2227 -104 2231 -84
rect 2295 -104 2299 -84
rect 2718 -102 2722 -82
rect 2786 -102 2790 -82
rect 3202 -4 3206 16
rect 2866 -104 2870 -84
rect 2934 -104 2938 -84
rect 3062 -100 3066 -80
rect 3130 -100 3134 -80
rect 3210 -102 3214 -82
rect 3278 -102 3282 -82
<< polycontact >>
rect 402 200 412 210
rect -86 122 -76 132
rect 258 124 268 134
rect 1385 202 1395 212
rect 624 128 634 138
rect 897 124 907 134
rect 1241 126 1251 136
rect 582 60 592 70
rect -136 -28 -126 -18
rect -60 -28 -50 -18
rect 472 6 482 16
rect 2407 204 2417 214
rect 1607 130 1617 140
rect 1919 126 1929 136
rect 2263 128 2273 138
rect 1565 62 1575 72
rect 208 -26 218 -16
rect 284 -26 294 -16
rect 847 -26 857 -16
rect 923 -26 933 -16
rect -128 -124 -118 -114
rect -26 -126 -16 -116
rect 1455 8 1465 18
rect 3390 206 3400 216
rect 2629 132 2639 142
rect 2902 128 2912 138
rect 3246 130 3256 140
rect 2587 64 2597 74
rect 1191 -24 1201 -14
rect 1267 -24 1277 -14
rect 216 -122 226 -112
rect 318 -124 328 -114
rect 1869 -24 1879 -14
rect 1945 -24 1955 -14
rect 855 -122 865 -112
rect 957 -124 967 -114
rect 2477 10 2487 20
rect 3612 134 3622 144
rect 3570 66 3580 76
rect 2213 -22 2223 -12
rect 2289 -22 2299 -12
rect 1199 -120 1209 -110
rect 1301 -122 1311 -112
rect 2852 -22 2862 -12
rect 2928 -22 2938 -12
rect 1877 -120 1887 -110
rect 1979 -122 1989 -112
rect 3460 12 3470 22
rect 3196 -20 3206 -10
rect 3272 -20 3282 -10
rect 2221 -118 2231 -108
rect 2323 -120 2333 -110
rect 2860 -118 2870 -108
rect 2962 -120 2972 -110
rect 3204 -116 3214 -106
rect 3306 -118 3316 -108
<< ndcontact >>
rect -286 112 -276 122
rect -194 112 -184 122
rect -100 106 -90 116
rect -66 106 -56 116
rect 58 114 68 124
rect 150 114 160 124
rect 244 108 254 118
rect 278 108 288 118
rect 697 114 707 124
rect 789 114 799 124
rect 394 38 404 48
rect 436 38 446 48
rect 486 38 496 48
rect 568 44 578 54
rect 602 44 612 54
rect -286 -42 -276 -32
rect -194 -42 -184 -32
rect -150 -44 -140 -34
rect -116 -44 -106 -34
rect 883 108 893 118
rect 917 108 927 118
rect 1041 116 1051 126
rect 1133 116 1143 126
rect 1227 110 1237 120
rect 1261 110 1271 120
rect 1719 116 1729 126
rect 1811 116 1821 126
rect 1377 40 1387 50
rect 1419 40 1429 50
rect 1469 40 1479 50
rect 1551 46 1561 56
rect 1585 46 1595 56
rect 58 -40 68 -30
rect 150 -40 160 -30
rect 194 -42 204 -32
rect 228 -42 238 -32
rect 697 -40 707 -30
rect 789 -40 799 -30
rect 833 -42 843 -32
rect 867 -42 877 -32
rect -286 -142 -276 -132
rect -244 -142 -234 -132
rect -194 -142 -184 -132
rect 1905 110 1915 120
rect 1939 110 1949 120
rect 2063 118 2073 128
rect 2155 118 2165 128
rect 2249 112 2259 122
rect 2283 112 2293 122
rect 2702 118 2712 128
rect 2794 118 2804 128
rect 2399 42 2409 52
rect 2441 42 2451 52
rect 2491 42 2501 52
rect 2573 48 2583 58
rect 2607 48 2617 58
rect 1041 -38 1051 -28
rect 1133 -38 1143 -28
rect 1177 -40 1187 -30
rect 1211 -40 1221 -30
rect -138 -144 -128 -134
rect -96 -144 -86 -134
rect -46 -144 -36 -134
rect 58 -140 68 -130
rect 100 -140 110 -130
rect 150 -140 160 -130
rect 1719 -38 1729 -28
rect 1811 -38 1821 -28
rect 1855 -40 1865 -30
rect 1889 -40 1899 -30
rect 206 -142 216 -132
rect 248 -142 258 -132
rect 298 -142 308 -132
rect 697 -140 707 -130
rect 739 -140 749 -130
rect 789 -140 799 -130
rect 2888 112 2898 122
rect 2922 112 2932 122
rect 3046 120 3056 130
rect 3138 120 3148 130
rect 3232 114 3242 124
rect 3266 114 3276 124
rect 3382 44 3392 54
rect 3424 44 3434 54
rect 3474 44 3484 54
rect 3556 50 3566 60
rect 3590 50 3600 60
rect 2063 -36 2073 -26
rect 2155 -36 2165 -26
rect 2199 -38 2209 -28
rect 2233 -38 2243 -28
rect 845 -142 855 -132
rect 887 -142 897 -132
rect 937 -142 947 -132
rect 1041 -138 1051 -128
rect 1083 -138 1093 -128
rect 1133 -138 1143 -128
rect 2702 -36 2712 -26
rect 2794 -36 2804 -26
rect 2838 -38 2848 -28
rect 2872 -38 2882 -28
rect 1189 -140 1199 -130
rect 1231 -140 1241 -130
rect 1281 -140 1291 -130
rect 1719 -138 1729 -128
rect 1761 -138 1771 -128
rect 1811 -138 1821 -128
rect 3046 -34 3056 -24
rect 3138 -34 3148 -24
rect 3182 -36 3192 -26
rect 3216 -36 3226 -26
rect 1867 -140 1877 -130
rect 1909 -140 1919 -130
rect 1959 -140 1969 -130
rect 2063 -136 2073 -126
rect 2105 -136 2115 -126
rect 2155 -136 2165 -126
rect 2211 -138 2221 -128
rect 2253 -138 2263 -128
rect 2303 -138 2313 -128
rect 2702 -136 2712 -126
rect 2744 -136 2754 -126
rect 2794 -136 2804 -126
rect 2850 -138 2860 -128
rect 2892 -138 2902 -128
rect 2942 -138 2952 -128
rect 3046 -134 3056 -124
rect 3088 -134 3098 -124
rect 3138 -134 3148 -124
rect 3194 -136 3204 -126
rect 3236 -136 3246 -126
rect 3286 -136 3296 -126
<< pdcontact >>
rect -286 150 -276 160
rect -244 150 -234 160
rect -194 150 -184 160
rect -100 144 -90 154
rect -66 144 -56 154
rect 58 152 68 162
rect 100 152 110 162
rect 150 152 160 162
rect 244 146 254 156
rect 278 146 288 156
rect -286 -4 -276 6
rect -244 -4 -234 6
rect 697 152 707 162
rect 739 152 749 162
rect 789 152 799 162
rect 883 146 893 156
rect 917 146 927 156
rect 1041 154 1051 164
rect 1083 154 1093 164
rect 1133 154 1143 164
rect 1227 148 1237 158
rect 1261 148 1271 158
rect 394 76 404 86
rect 486 76 496 86
rect 568 82 578 92
rect 602 82 612 92
rect -194 -4 -184 6
rect -150 -6 -140 4
rect -116 -6 -106 4
rect 58 -2 68 8
rect 100 -2 110 8
rect 150 -2 160 8
rect 194 -4 204 6
rect -286 -104 -276 -94
rect 228 -4 238 6
rect 697 -2 707 8
rect 739 -2 749 8
rect 1719 154 1729 164
rect 1761 154 1771 164
rect 1811 154 1821 164
rect 1905 148 1915 158
rect 1939 148 1949 158
rect 2063 156 2073 166
rect 2105 156 2115 166
rect 2155 156 2165 166
rect 2249 150 2259 160
rect 2283 150 2293 160
rect 1377 78 1387 88
rect 1469 78 1479 88
rect 1551 84 1561 94
rect 1585 84 1595 94
rect 789 -2 799 8
rect 833 -4 843 6
rect -194 -104 -184 -94
rect -138 -106 -128 -96
rect -46 -106 -36 -96
rect 58 -102 68 -92
rect 867 -4 877 6
rect 1041 0 1051 10
rect 1083 0 1093 10
rect 1133 0 1143 10
rect 1177 -2 1187 8
rect 150 -102 160 -92
rect 206 -104 216 -94
rect 298 -104 308 -94
rect 697 -102 707 -92
rect 1211 -2 1221 8
rect 1719 0 1729 10
rect 1761 0 1771 10
rect 2702 156 2712 166
rect 2744 156 2754 166
rect 2794 156 2804 166
rect 2888 150 2898 160
rect 2922 150 2932 160
rect 3046 158 3056 168
rect 3088 158 3098 168
rect 3138 158 3148 168
rect 3232 152 3242 162
rect 3266 152 3276 162
rect 2399 80 2409 90
rect 2491 80 2501 90
rect 2573 86 2583 96
rect 2607 86 2617 96
rect 1811 0 1821 10
rect 1855 -2 1865 8
rect 789 -102 799 -92
rect 845 -104 855 -94
rect 937 -104 947 -94
rect 1041 -100 1051 -90
rect 1889 -2 1899 8
rect 2063 2 2073 12
rect 2105 2 2115 12
rect 2155 2 2165 12
rect 2199 0 2209 10
rect 1133 -100 1143 -90
rect 1189 -102 1199 -92
rect 1281 -102 1291 -92
rect 1719 -100 1729 -90
rect 2233 0 2243 10
rect 2702 2 2712 12
rect 2744 2 2754 12
rect 3382 82 3392 92
rect 3474 82 3484 92
rect 3556 88 3566 98
rect 3590 88 3600 98
rect 2794 2 2804 12
rect 2838 0 2848 10
rect 1811 -100 1821 -90
rect 1867 -102 1877 -92
rect 1959 -102 1969 -92
rect 2063 -98 2073 -88
rect 2872 0 2882 10
rect 3046 4 3056 14
rect 3088 4 3098 14
rect 3138 4 3148 14
rect 3182 2 3192 12
rect 2155 -98 2165 -88
rect 2211 -100 2221 -90
rect 2303 -100 2313 -90
rect 2702 -98 2712 -88
rect 3216 2 3226 12
rect 2794 -98 2804 -88
rect 2850 -100 2860 -90
rect 2942 -100 2952 -90
rect 3046 -96 3056 -86
rect 3138 -96 3148 -86
rect 3194 -98 3204 -88
rect 3286 -98 3296 -88
<< m2contact >>
rect 326 200 336 210
rect 1309 202 1319 212
rect 2331 204 2341 214
rect 3314 206 3324 216
rect -48 122 -38 132
rect 296 124 306 134
rect 320 94 330 104
rect 382 94 392 104
rect 935 124 945 134
rect 444 6 454 16
rect 1279 126 1289 136
rect 1303 96 1313 106
rect 1365 96 1375 106
rect 1957 126 1967 136
rect 1427 8 1437 18
rect 2301 128 2311 138
rect 2325 98 2335 108
rect 2387 98 2397 108
rect 2940 128 2950 138
rect 2449 10 2459 20
rect 3284 130 3294 140
rect 3308 100 3318 110
rect 3370 100 3380 110
rect 3432 12 3442 22
<< labels >>
rlabel metal1 -305 101 -305 101 3 gnd
rlabel metal1 -291 173 -291 173 1 vdd
rlabel polysilicon 144 224 144 224 5 cin
rlabel polysilicon 715 226 715 226 1 a2
rlabel polysilicon 783 227 783 227 1 b2
rlabel polysilicon -267 223 -267 223 1 a1
rlabel polysilicon -200 222 -200 222 1 b1
rlabel polysilicon 3618 166 3618 166 7 cout
rlabel polysilicon 1737 227 1737 227 1 a3
rlabel polysilicon 1805 229 1805 229 1 b3
rlabel polysilicon 2720 228 2720 228 1 a4
rlabel polysilicon 2788 229 2788 229 1 b4
rlabel polysilicon 3327 -112 3327 -112 1 s4
rlabel polysilicon 2344 -114 2344 -114 1 s3
rlabel polysilicon 1322 -116 1322 -116 1 s2
rlabel polysilicon 338 -118 338 -118 1 s1
<< end >>
